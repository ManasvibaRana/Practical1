<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-17.8,-91.2333,176.6,-189.5</PageViewport>
<gate>
<ID>2</ID>
<type>AA_MUX_2x1</type>
<position>25,-18.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>3 </output>
<input>
<ID>SEL_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>53,-18.5</position>
<gparam>LABEL_TEXT 1 * 4 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>HA_JUNC_2</type>
<position>-27.5,-24.5</position>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>67.5,-9.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>15,-17</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>75.5,-9.5</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>15,-20</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>75.5,-6.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>32,-18.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>67.5,-6.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>25,-10.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>11.5,-20</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>11.5,-16.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>25,-7.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>0,-18</position>
<gparam>LABEL_TEXT 2 * 1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>-0.5,-35</position>
<gparam>LABEL_TEXT 4 * 1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AE_MUX_4x1</type>
<position>24,-36</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>8 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>6 </input>
<output>
<ID>OUT</ID>12 </output>
<input>
<ID>SEL_0</ID>11 </input>
<input>
<ID>SEL_1</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>13.5,-31</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>13.5,-34</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>13.5,-37.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>13.5,-41</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>24,-24</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>27,-24</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_AND3</type>
<position>90.5,-16.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>31 </input>
<input>
<ID>IN_2</ID>4 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>32.5,-36</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>10,-40.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>10,-37</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>10,-30.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>10,-33.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>29,-44</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>26.5,-44</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>-1,-55.5</position>
<gparam>LABEL_TEXT 8 * 1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND3</type>
<position>90.5,-25</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<input>
<ID>IN_2</ID>4 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>39</ID>
<type>AI_MUX_8x1</type>
<position>27.5,-62.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>20 </input>
<input>
<ID>IN_2</ID>19 </input>
<input>
<ID>IN_3</ID>22 </input>
<input>
<ID>IN_4</ID>17 </input>
<input>
<ID>IN_5</ID>16 </input>
<input>
<ID>IN_6</ID>14 </input>
<input>
<ID>IN_7</ID>13 </input>
<output>
<ID>OUT</ID>26 </output>
<input>
<ID>SEL_0</ID>23 </input>
<input>
<ID>SEL_1</ID>24 </input>
<input>
<ID>SEL_2</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>12.5,-53.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_TOGGLE</type>
<position>12.5,-56</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>12.5,-58.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>12.5,-61</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>12.5,-63.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>12.5,-66</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>12.5,-68.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>12.5,-71</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>28.5,-46.5</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>26.5,-46.5</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>24.5,-46.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>51</ID>
<type>GA_LED</type>
<position>35,-62.5</position>
<input>
<ID>N_in0</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>27,-21.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>24,-21.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>24,-44</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>9,-71</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>9,-68.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>9,-66</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>9,-63.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>9,-61</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>9,-58.5</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>9,-56</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>9,-53.5</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_AND3</type>
<position>91,-33.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>30 </input>
<input>
<ID>IN_2</ID>4 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_AND3</type>
<position>91,-43</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>32 </input>
<input>
<ID>IN_2</ID>4 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_TOGGLE</type>
<position>83.5,-9.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>83.5,-6.5</position>
<gparam>LABEL_TEXT Din</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>68</ID>
<type>AE_SMALL_INVERTER</type>
<position>71,-13</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>70</ID>
<type>AE_SMALL_INVERTER</type>
<position>79,-13</position>
<input>
<ID>IN_0</ID>32 </input>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>72</ID>
<type>GA_LED</type>
<position>98,-16.5</position>
<input>
<ID>N_in0</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>GA_LED</type>
<position>97.5,-25</position>
<input>
<ID>N_in0</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>GA_LED</type>
<position>97.5,-33.5</position>
<input>
<ID>N_in0</ID>34 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>GA_LED</type>
<position>98,-43</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>102,-16.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>101.5,-25</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>101,-33</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>101,-42.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>52.5,-70</position>
<gparam>LABEL_TEXT 1 * 8 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>66.5,-57</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_TOGGLE</type>
<position>74.5,-57</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>82,-57</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_TOGGLE</type>
<position>89.5,-57</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>89.5,-54</position>
<gparam>LABEL_TEXT Din</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>74.5,-54</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>82,-54.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>66.5,-54</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_AND4</type>
<position>102,-65.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>54 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>37 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_AND4</type>
<position>102,-74.5</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>54 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>37 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_AND4</type>
<position>102,-83.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>57 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>37 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_AND4</type>
<position>102,-92.5</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>57 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>37 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_AND4</type>
<position>102,-101.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>54 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>37 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_AND4</type>
<position>102,-110.5</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>54 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>37 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_AND4</type>
<position>102.5,-119.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>57 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>37 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_AND4</type>
<position>102,-128.5</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>57 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>37 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>109</ID>
<type>GA_LED</type>
<position>110.5,-65.5</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>GA_LED</type>
<position>110,-74.5</position>
<input>
<ID>N_in0</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>GA_LED</type>
<position>110,-83.5</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>GA_LED</type>
<position>110,-92.5</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>GA_LED</type>
<position>110,-101.5</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>GA_LED</type>
<position>110.5,-110.5</position>
<input>
<ID>N_in0</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>GA_LED</type>
<position>110.5,-119.5</position>
<input>
<ID>N_in0</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>GA_LED</type>
<position>110.5,-128.5</position>
<input>
<ID>N_in0</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AE_SMALL_INVERTER</type>
<position>85,-61</position>
<input>
<ID>IN_0</ID>56 </input>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_SMALL_INVERTER</type>
<position>78.5,-61</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>120</ID>
<type>AE_SMALL_INVERTER</type>
<position>70.5,-61</position>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>114,-65</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>113.5,-74</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>2,-168.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_LABEL</type>
<position>2,-165</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>125</ID>
<type>AA_LABEL</type>
<position>113.5,-101.5</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>114,-110</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>114,-119</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>114.5,-128</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_LABEL</type>
<position>-1.5,-141</position>
<gparam>LABEL_TEXT 4 * 1 using 2*1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_MUX_2x1</type>
<position>14,-154.5</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>70 </output>
<input>
<ID>SEL_0</ID>64 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_MUX_2x1</type>
<position>13.5,-166.5</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>71 </output>
<input>
<ID>SEL_0</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_MUX_2x1</type>
<position>24,-160</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>71 </input>
<output>
<ID>OUT</ID>73 </output>
<input>
<ID>SEL_0</ID>72 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_TOGGLE</type>
<position>5,-153</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_TOGGLE</type>
<position>5,-156</position>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_TOGGLE</type>
<position>5.5,-165.5</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_TOGGLE</type>
<position>5.5,-168.5</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_TOGGLE</type>
<position>14,-147</position>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>146</ID>
<type>AA_TOGGLE</type>
<position>13.5,-160</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_TOGGLE</type>
<position>24,-153.5</position>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>149</ID>
<type>GA_LED</type>
<position>28.5,-160</position>
<input>
<ID>N_in0</ID>73 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>AA_LABEL</type>
<position>2,-156</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>151</ID>
<type>AA_LABEL</type>
<position>2,-152</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>152</ID>
<type>AA_LABEL</type>
<position>14,-144.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>13.5,-157.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>154</ID>
<type>AA_LABEL</type>
<position>24,-150</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-17.5,23,-17.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>17 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>17,-17.5,17,-17</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-19.5,23,-19.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>17 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>17,-20,17,-19.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-18.5,31,-18.5</points>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-45,83.5,-11.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>-45 5</intersection>
<intersection>-35.5 6</intersection>
<intersection>-27 7</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-18.5,87.5,-18.5</points>
<connection>
<GID>29</GID>
<name>IN_2</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>83.5,-45,88,-45</points>
<connection>
<GID>64</GID>
<name>IN_2</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>83.5,-35.5,88,-35.5</points>
<connection>
<GID>63</GID>
<name>IN_2</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>83.5,-27,87.5,-27</points>
<connection>
<GID>38</GID>
<name>IN_2</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-16,25,-12.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-33,18,-31</points>
<intersection>-33 1</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-33,21,-33</points>
<connection>
<GID>21</GID>
<name>IN_3</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-31,18,-31</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-35,18,-34</points>
<intersection>-35 1</intersection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-35,21,-35</points>
<connection>
<GID>21</GID>
<name>IN_2</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-34,18,-34</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-37.5,18,-37</points>
<intersection>-37.5 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-37,21,-37</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-37.5,18,-37.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-41,18,-39</points>
<intersection>-41 1</intersection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,-41,18,-41</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-39,21,-39</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-31,24,-26</points>
<connection>
<GID>21</GID>
<name>SEL_1</name></connection>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-31,25,-28.5</points>
<connection>
<GID>21</GID>
<name>SEL_0</name></connection>
<intersection>-28.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>27,-28.5,27,-26</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>25,-28.5,27,-28.5</points>
<intersection>25 0</intersection>
<intersection>27 1</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-36,31.5,-36</points>
<connection>
<GID>30</GID>
<name>N_in0</name></connection>
<connection>
<GID>21</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-59,23,-53.5</points>
<intersection>-59 1</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-59,24.5,-59</points>
<connection>
<GID>39</GID>
<name>IN_7</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-53.5,23,-53.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14.5,-56,22,-56</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>22 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>22,-60,22,-56</points>
<intersection>-60 10</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>22,-60,24.5,-60</points>
<connection>
<GID>39</GID>
<name>IN_6</name></connection>
<intersection>22 9</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-61,19.5,-58</points>
<intersection>-61 1</intersection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-61,24.5,-61</points>
<connection>
<GID>39</GID>
<name>IN_5</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-58,19.5,-58</points>
<intersection>14.5 3</intersection>
<intersection>19.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14.5,-58.5,14.5,-58</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>-58 2</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-62,18.5,-61</points>
<intersection>-62 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-61,18.5,-61</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-62,24.5,-62</points>
<connection>
<GID>39</GID>
<name>IN_4</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-66,17,-64</points>
<intersection>-66 1</intersection>
<intersection>-64 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-66,17,-66</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-64,24.5,-64</points>
<connection>
<GID>39</GID>
<name>IN_2</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-68.5,18,-65</points>
<intersection>-68.5 1</intersection>
<intersection>-65 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-68.5,18,-68.5</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-65,24.5,-65</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-71,19.5,-66</points>
<intersection>-71 1</intersection>
<intersection>-66 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-71,19.5,-71</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-66,24.5,-66</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-63.5,19.5,-63</points>
<intersection>-63.5 1</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-63.5,19.5,-63.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-63,24.5,-63</points>
<connection>
<GID>39</GID>
<name>IN_3</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-57,28.5,-48.5</points>
<connection>
<GID>39</GID>
<name>SEL_0</name></connection>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-57,27.5,-53.5</points>
<connection>
<GID>39</GID>
<name>SEL_1</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>26.5,-53.5,26.5,-48.5</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-53.5,27.5,-53.5</points>
<intersection>26.5 1</intersection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-57,25.5,-52.5</points>
<intersection>-57 3</intersection>
<intersection>-52.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>24.5,-52.5,24.5,-48.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>-52.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-52.5,25.5,-52.5</points>
<intersection>24.5 1</intersection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25.5,-57,26.5,-57</points>
<connection>
<GID>39</GID>
<name>SEL_2</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-62.5,34,-62.5</points>
<connection>
<GID>51</GID>
<name>N_in0</name></connection>
<connection>
<GID>39</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-41,67.5,-11.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>-41 3</intersection>
<intersection>-31.5 1</intersection>
<intersection>-13 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-31.5,88,-31.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>67.5,-41,88,-41</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>67.5,-13,69,-13</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,-16.5,97,-16.5</points>
<connection>
<GID>72</GID>
<name>N_in0</name></connection>
<connection>
<GID>29</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-14.5,84,-13</points>
<intersection>-14.5 1</intersection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,-14.5,87.5,-14.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>81.5 3</intersection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81,-13,84,-13</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>84 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>81.5,-33.5,81.5,-14.5</points>
<intersection>-33.5 4</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>81.5,-33.5,88,-33.5</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>81.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-23,73,-13</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>-23 3</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-16.5,87.5,-16.5</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>73,-23,87.5,-23</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-43,75.5,-11.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-43 5</intersection>
<intersection>-25 3</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-13,77,-13</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>75.5,-25,87.5,-25</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>75.5,-43,88,-43</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,-25,96.5,-25</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<connection>
<GID>73</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-33.5,96.5,-33.5</points>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<connection>
<GID>74</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-43,97,-43</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<connection>
<GID>75</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-131.5,89.5,-59</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<intersection>-131.5 9</intersection>
<intersection>-122.5 8</intersection>
<intersection>-113.5 7</intersection>
<intersection>-104.5 6</intersection>
<intersection>-95.5 5</intersection>
<intersection>-86.5 4</intersection>
<intersection>-77.5 3</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-68.5,99,-68.5</points>
<connection>
<GID>100</GID>
<name>IN_3</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>89.5,-77.5,99,-77.5</points>
<connection>
<GID>101</GID>
<name>IN_3</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>89.5,-86.5,99,-86.5</points>
<connection>
<GID>102</GID>
<name>IN_3</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>89.5,-95.5,99,-95.5</points>
<connection>
<GID>103</GID>
<name>IN_3</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>89.5,-104.5,99,-104.5</points>
<connection>
<GID>104</GID>
<name>IN_3</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>89.5,-113.5,99,-113.5</points>
<connection>
<GID>105</GID>
<name>IN_3</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>89.5,-122.5,99.5,-122.5</points>
<connection>
<GID>106</GID>
<name>IN_3</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>89.5,-131.5,99,-131.5</points>
<connection>
<GID>107</GID>
<name>IN_3</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-65.5,109.5,-65.5</points>
<connection>
<GID>109</GID>
<name>N_in0</name></connection>
<connection>
<GID>100</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-74.5,109,-74.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<connection>
<GID>110</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-83.5,109,-83.5</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<connection>
<GID>111</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-92.5,109,-92.5</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<connection>
<GID>112</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-101.5,109,-101.5</points>
<connection>
<GID>104</GID>
<name>OUT</name></connection>
<connection>
<GID>113</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-110.5,109.5,-110.5</points>
<connection>
<GID>105</GID>
<name>OUT</name></connection>
<connection>
<GID>114</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105.5,-119.5,109.5,-119.5</points>
<connection>
<GID>115</GID>
<name>N_in0</name></connection>
<connection>
<GID>106</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-128.5,109.5,-128.5</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<connection>
<GID>116</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80.5,-64.5,99,-64.5</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>80.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>80.5,-109.5,80.5,-61</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 9</intersection>
<intersection>-100.5 7</intersection>
<intersection>-73.5 5</intersection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>80.5,-73.5,99,-73.5</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>80.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>80.5,-100.5,99,-100.5</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<intersection>80.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>80.5,-109.5,99,-109.5</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>80.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-93.5,72.5,-61</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<intersection>-93.5 8</intersection>
<intersection>-84.5 6</intersection>
<intersection>-75.5 4</intersection>
<intersection>-66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-66.5,99,-66.5</points>
<connection>
<GID>100</GID>
<name>IN_2</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>72.5,-75.5,99,-75.5</points>
<connection>
<GID>101</GID>
<name>IN_2</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>72.5,-84.5,99,-84.5</points>
<connection>
<GID>102</GID>
<name>IN_2</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>72.5,-93.5,99,-93.5</points>
<connection>
<GID>103</GID>
<name>IN_2</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-125.5,82,-59</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>-125.5 9</intersection>
<intersection>-107.5 5</intersection>
<intersection>-89.5 3</intersection>
<intersection>-71.5 1</intersection>
<intersection>-61 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-71.5,99,-71.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>82,-89.5,99,-89.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>82,-107.5,99,-107.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>82,-61,83,-61</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>82,-125.5,99,-125.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-127.5,74.5,-59</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>-127.5 5</intersection>
<intersection>-118.5 7</intersection>
<intersection>-91.5 3</intersection>
<intersection>-82.5 1</intersection>
<intersection>-61 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-82.5,99,-82.5</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>74.5,-91.5,99,-91.5</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>74.5,-127.5,99,-127.5</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>74.5,-118.5,99.5,-118.5</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>74.5,-61,76.5,-61</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-129.5,66.5,-59</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>-129.5 7</intersection>
<intersection>-120.5 5</intersection>
<intersection>-111.5 3</intersection>
<intersection>-102.5 1</intersection>
<intersection>-61 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-102.5,99,-102.5</points>
<connection>
<GID>104</GID>
<name>IN_2</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>66.5,-111.5,99,-111.5</points>
<connection>
<GID>105</GID>
<name>IN_2</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>66.5,-120.5,99.5,-120.5</points>
<connection>
<GID>106</GID>
<name>IN_2</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>66.5,-129.5,99,-129.5</points>
<connection>
<GID>107</GID>
<name>IN_2</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>66.5,-61,68.5,-61</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87,-62.5,99,-62.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>87 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>87,-116.5,87,-61</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>-116.5 9</intersection>
<intersection>-98.5 7</intersection>
<intersection>-80.5 5</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>87,-80.5,99,-80.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>87 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>87,-98.5,99,-98.5</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>87 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>87,-116.5,99.5,-116.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>87 3</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-153.5,9.5,-153</points>
<intersection>-153.5 1</intersection>
<intersection>-153 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,-153.5,12,-153.5</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-153,9.5,-153</points>
<connection>
<GID>138</GID>
<name>OUT_0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-156,9.5,-155.5</points>
<intersection>-156 2</intersection>
<intersection>-155.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,-155.5,12,-155.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-156,9.5,-156</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-165.5,11.5,-165.5</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-168.5,9.5,-167.5</points>
<intersection>-168.5 1</intersection>
<intersection>-167.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,-168.5,9.5,-168.5</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-167.5,11.5,-167.5</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-152,14,-149</points>
<connection>
<GID>145</GID>
<name>OUT_0</name></connection>
<intersection>-152 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>14,-152,14,-152</points>
<connection>
<GID>132</GID>
<name>SEL_0</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-164,13.5,-162</points>
<connection>
<GID>146</GID>
<name>OUT_0</name></connection>
<intersection>-164 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>13.5,-164,13.5,-164</points>
<connection>
<GID>134</GID>
<name>SEL_0</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-161,19,-154.5</points>
<intersection>-161 1</intersection>
<intersection>-154.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-161,22,-161</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-154.5,19,-154.5</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-166.5,18.5,-159</points>
<intersection>-166.5 2</intersection>
<intersection>-159 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-159,22,-159</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-166.5,18.5,-166.5</points>
<connection>
<GID>134</GID>
<name>OUT</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-157.5,24,-155.5</points>
<connection>
<GID>136</GID>
<name>SEL_0</name></connection>
<connection>
<GID>147</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-160,27.5,-160</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<connection>
<GID>149</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,2.29719e-006,145.8,-73.7</PageViewport></page 1>
<page 2>
<PageViewport>0,2.29719e-006,145.8,-73.7</PageViewport></page 2>
<page 3>
<PageViewport>0,2.29719e-006,145.8,-73.7</PageViewport></page 3>
<page 4>
<PageViewport>0,2.29719e-006,145.8,-73.7</PageViewport></page 4>
<page 5>
<PageViewport>0,2.29719e-006,145.8,-73.7</PageViewport></page 5>
<page 6>
<PageViewport>0,2.29719e-006,145.8,-73.7</PageViewport></page 6>
<page 7>
<PageViewport>0,2.29719e-006,145.8,-73.7</PageViewport></page 7>
<page 8>
<PageViewport>0,2.29719e-006,145.8,-73.7</PageViewport></page 8>
<page 9>
<PageViewport>0,2.29719e-006,145.8,-73.7</PageViewport></page 9></circuit>