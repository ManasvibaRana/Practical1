<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-39.4735,-403.898,154.926,-502.164</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>-26,42</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>-43,45</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>-43,39</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>-20,41.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>-43,29.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>-44,8.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>3,-16.5</position>
<gparam>LABEL_TEXT NAND AS A UNIVERSAL GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>-50,45.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>-50,39.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>-43,24</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>23</ID>
<type>AE_OR2</type>
<position>-26.5,26.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>-44,13.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>-19.5,26.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>-51,30</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>-50.5,24</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>-37.5,35</position>
<gparam>LABEL_TEXT OR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>-36,19.5</position>
<gparam>LABEL_TEXT NAND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>-10,42</position>
<gparam>LABEL_TEXT Y = A*B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>-8.5,26.5</position>
<gparam>LABEL_TEXT Y = A+B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>BA_NAND2</type>
<position>-26.5,11.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>-20,11.5</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>-5.5,16</position>
<gparam>LABEL_TEXT ____</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>-8.5,12.5</position>
<gparam>LABEL_TEXT Y = A*B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>-51.5,14</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>-51.5,9</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>-36.5,3</position>
<gparam>LABEL_TEXT NOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>-44,-3</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>-44,-9</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>BE_NOR2</type>
<position>-26.5,-6</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>GA_LED</type>
<position>-21,-6</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>-51.5,-2.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>-51.5,-8.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>-10.5,-5.5</position>
<gparam>LABEL_TEXT Y = A+B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>-8,-2.5</position>
<gparam>LABEL_TEXT ____</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>18,45.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_TOGGLE</type>
<position>18,40.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>61</ID>
<type>GA_LED</type>
<position>47.5,43.5</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AO_XNOR2</type>
<position>38.5,43.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>30.5,51.5</position>
<gparam>LABEL_TEXT XOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>10,46</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>10,41</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>58.5,44</position>
<gparam>LABEL_TEXT Y = AB + AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>56.5,47</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>66.5,47</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>30,34</position>
<gparam>LABEL_TEXT XNOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>72</ID>
<type>BA_NAND2</type>
<position>-1,-32</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>-12,-32</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>76</ID>
<type>GA_LED</type>
<position>7,-32</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>-35,-30.5</position>
<gparam>LABEL_TEXT NAND AS A NOT GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>79</ID>
<type>BA_NAND2</type>
<position>-1,-41.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_TOGGLE</type>
<position>-12,-40</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_TOGGLE</type>
<position>-12,-44</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>84</ID>
<type>BA_NAND2</type>
<position>10,-41.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>GA_LED</type>
<position>17.5,-41.5</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>-34,-42</position>
<gparam>LABEL_TEXT NAND AS A AND GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>87</ID>
<type>BA_NAND2</type>
<position>-1.5,-51.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>88</ID>
<type>BA_NAND2</type>
<position>-1.5,-59</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_TOGGLE</type>
<position>-12,-51.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_TOGGLE</type>
<position>-12,-59</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>91</ID>
<type>BA_NAND2</type>
<position>9,-55</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>GA_LED</type>
<position>17,-55</position>
<input>
<ID>N_in0</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_LABEL</type>
<position>-34,-55</position>
<gparam>LABEL_TEXT NAND AS A OR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>94</ID>
<type>BA_NAND2</type>
<position>-1,-68</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>BA_NAND2</type>
<position>-1,-76.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>96</ID>
<type>BA_NAND2</type>
<position>9.5,-71.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>97</ID>
<type>BA_NAND2</type>
<position>19,-71.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_TOGGLE</type>
<position>-12,-68</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_TOGGLE</type>
<position>-12,-76.5</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>100</ID>
<type>GA_LED</type>
<position>27.5,-71.5</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>AA_LABEL</type>
<position>-33,-72</position>
<gparam>LABEL_TEXT NAND AS A NOR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>110</ID>
<type>AA_TOGGLE</type>
<position>-12,-85.5</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_TOGGLE</type>
<position>-12,-93.5</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>112</ID>
<type>BA_NAND2</type>
<position>-2,-89.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>BA_NAND2</type>
<position>7.5,-86</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>BA_NAND2</type>
<position>8,-92.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>BA_NAND2</type>
<position>17.5,-89</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>GA_LED</type>
<position>26.5,-89</position>
<input>
<ID>N_in0</ID>50 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>-33.5,-89.5</position>
<gparam>LABEL_TEXT NAND AS A XOR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_TOGGLE</type>
<position>-12,-102</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_TOGGLE</type>
<position>-12,-110</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>120</ID>
<type>BA_NAND2</type>
<position>-2,-106</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>BA_NAND2</type>
<position>7.5,-102.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>BA_NAND2</type>
<position>8,-109</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>BA_NAND2</type>
<position>17.5,-105.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>GA_LED</type>
<position>33.5,-105.5</position>
<input>
<ID>N_in0</ID>58 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>BA_NAND2</type>
<position>26,-105.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>-32.5,-105</position>
<gparam>LABEL_TEXT NAND AS A XNOR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>-8.5,-121.5</position>
<gparam>LABEL_TEXT NOR AS A UNIVERSAL GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>-34,-137</position>
<gparam>LABEL_TEXT NOR AS A NOT GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>130</ID>
<type>BE_NOR2</type>
<position>-1.5,-137.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>131</ID>
<type>AA_TOGGLE</type>
<position>-12.5,-137.5</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>133</ID>
<type>GA_LED</type>
<position>3.5,-137.5</position>
<input>
<ID>N_in0</ID>60 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>BE_NOR2</type>
<position>-2,-147.5</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_TOGGLE</type>
<position>-12.5,-145.5</position>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>137</ID>
<type>AA_TOGGLE</type>
<position>-12.5,-150</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>140</ID>
<type>BE_NOR2</type>
<position>7,-147.5</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>141</ID>
<type>GA_LED</type>
<position>13,-147.5</position>
<input>
<ID>N_in0</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>AA_LABEL</type>
<position>-33,-147.5</position>
<gparam>LABEL_TEXT NOR AS A OR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>144</ID>
<type>BE_NOR2</type>
<position>-3,-159</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_TOGGLE</type>
<position>-13,-159</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>146</ID>
<type>BE_NOR2</type>
<position>-3,-166</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_TOGGLE</type>
<position>-13,-166</position>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>148</ID>
<type>BE_NOR2</type>
<position>6.5,-162.5</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>149</ID>
<type>GA_LED</type>
<position>13.5,-162.5</position>
<input>
<ID>N_in0</ID>68 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>AA_LABEL</type>
<position>-33,-162.5</position>
<gparam>LABEL_TEXT NOR AS A AND GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>151</ID>
<type>BE_NOR2</type>
<position>-3,-176.5</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>152</ID>
<type>AA_TOGGLE</type>
<position>-13,-176.5</position>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>153</ID>
<type>BE_NOR2</type>
<position>-3,-183.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>73 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>154</ID>
<type>AA_TOGGLE</type>
<position>-13,-183.5</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>155</ID>
<type>BE_NOR2</type>
<position>6.5,-180</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>BE_NOR2</type>
<position>15.5,-180</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>GA_LED</type>
<position>21.5,-180</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>AA_LABEL</type>
<position>-32.5,-180</position>
<gparam>LABEL_TEXT NOR AS A NAND GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>160</ID>
<type>BE_NOR2</type>
<position>-4,-198.5</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>BE_NOR2</type>
<position>4,-193</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>162</ID>
<type>BE_NOR2</type>
<position>4,-204</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>163</ID>
<type>AA_TOGGLE</type>
<position>-14.5,-194.5</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>164</ID>
<type>AA_TOGGLE</type>
<position>-14.5,-203</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>165</ID>
<type>BE_NOR2</type>
<position>13.5,-198</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>166</ID>
<type>BE_NOR2</type>
<position>22.5,-198</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>167</ID>
<type>GA_LED</type>
<position>27.5,-198</position>
<input>
<ID>N_in0</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AA_LABEL</type>
<position>-34.5,-198.5</position>
<gparam>LABEL_TEXT NOR AS A XOR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>169</ID>
<type>BE_NOR2</type>
<position>-4,-219.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>BE_NOR2</type>
<position>4,-214</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>BE_NOR2</type>
<position>4,-225</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_TOGGLE</type>
<position>-15.5,-215</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_TOGGLE</type>
<position>-16.5,-223.5</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>174</ID>
<type>BE_NOR2</type>
<position>13.5,-219</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>GA_LED</type>
<position>21.5,-219</position>
<input>
<ID>N_in0</ID>93 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>AA_LABEL</type>
<position>-35,-219</position>
<gparam>LABEL_TEXT NOR AS A XNOR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>179</ID>
<type>AA_LABEL</type>
<position>1.5,-237.5</position>
<gparam>LABEL_TEXT HALF ADDER</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>181</ID>
<type>AO_XNOR2</type>
<position>-4,-250.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_TOGGLE</type>
<position>-14.5,-248</position>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>183</ID>
<type>AA_TOGGLE</type>
<position>-14.5,-253.5</position>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>184</ID>
<type>GA_LED</type>
<position>4,-250.5</position>
<input>
<ID>N_in0</ID>96 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>-24,-247.5</position>
<gparam>LABEL_TEXT INPUT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>AA_LABEL</type>
<position>-24,-253.5</position>
<gparam>LABEL_TEXT INPUT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>188</ID>
<type>AA_LABEL</type>
<position>17.5,-250</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>189</ID>
<type>AA_LABEL</type>
<position>20.5,-250.5</position>
<gparam>LABEL_TEXT SUM = AB + AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>191</ID>
<type>AA_LABEL</type>
<position>21,-247.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>192</ID>
<type>AA_LABEL</type>
<position>31,-247.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>194</ID>
<type>AA_LABEL</type>
<position>0,-264.5</position>
<gparam>LABEL_TEXT AOI IMPLIMENTATION</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>196</ID>
<type>AA_TOGGLE</type>
<position>-27.5,-271</position>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_AND2</type>
<position>-4.5,-257.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>GA_LED</type>
<position>3.5,-257.5</position>
<input>
<ID>N_in0</ID>98 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>AA_LABEL</type>
<position>18,-257</position>
<gparam>LABEL_TEXT CARRY = AB </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>AA_TOGGLE</type>
<position>-16,-271</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>206</ID>
<type>AE_SMALL_INVERTER</type>
<position>-24.5,-275.5</position>
<input>
<ID>IN_0</ID>104 </input>
<output>
<ID>OUT_0</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>207</ID>
<type>AE_SMALL_INVERTER</type>
<position>-13,-274.5</position>
<input>
<ID>IN_0</ID>103 </input>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_LABEL</type>
<position>-27.5,-267.5</position>
<gparam>LABEL_TEXT INPUT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AA_LABEL</type>
<position>-15,-267.5</position>
<gparam>LABEL_TEXT INPUT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>AA_AND2</type>
<position>1.5,-280</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>AA_AND2</type>
<position>1.5,-287.5</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>AE_OR2</type>
<position>13.5,-283</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>107 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>217</ID>
<type>GA_LED</type>
<position>21.5,-283</position>
<input>
<ID>N_in0</ID>108 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_AND2</type>
<position>0.5,-298</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>221</ID>
<type>GA_LED</type>
<position>13,-298</position>
<input>
<ID>N_in0</ID>112 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>34.5,-282</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>AA_LABEL</type>
<position>37.5,-282.5</position>
<gparam>LABEL_TEXT SUM = AB + AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>226</ID>
<type>AA_LABEL</type>
<position>37.5,-279.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>227</ID>
<type>AA_LABEL</type>
<position>48,-279.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>228</ID>
<type>AA_LABEL</type>
<position>0.5,-305</position>
<gparam>LABEL_TEXT NAND IMPLIMENTATION</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>229</ID>
<type>AA_TOGGLE</type>
<position>-27.5,-312.5</position>
<output>
<ID>OUT_0</ID>113 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>231</ID>
<type>AA_TOGGLE</type>
<position>-13.5,-312.5</position>
<output>
<ID>OUT_0</ID>115 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>233</ID>
<type>BA_NAND2</type>
<position>-21,-317</position>
<input>
<ID>IN_0</ID>113 </input>
<input>
<ID>IN_1</ID>113 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>235</ID>
<type>BA_NAND2</type>
<position>-8,-317.5</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>236</ID>
<type>BA_NAND2</type>
<position>3,-325</position>
<input>
<ID>IN_0</ID>113 </input>
<input>
<ID>IN_1</ID>114 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>BA_NAND2</type>
<position>3.5,-333.5</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>116 </input>
<output>
<ID>OUT</ID>118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>238</ID>
<type>BA_NAND2</type>
<position>15,-329</position>
<input>
<ID>IN_0</ID>117 </input>
<input>
<ID>IN_1</ID>118 </input>
<output>
<ID>OUT</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>239</ID>
<type>GA_LED</type>
<position>23,-329</position>
<input>
<ID>N_in0</ID>119 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>240</ID>
<type>AA_LABEL</type>
<position>36,-328</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>241</ID>
<type>AA_LABEL</type>
<position>39,-328.5</position>
<gparam>LABEL_TEXT SUM = AB + AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>AA_LABEL</type>
<position>39.5,-325.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>243</ID>
<type>AA_LABEL</type>
<position>49.5,-325.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>BA_NAND2</type>
<position>4,-344</position>
<input>
<ID>IN_0</ID>113 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>247</ID>
<type>BA_NAND2</type>
<position>18.5,-344</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>120 </input>
<output>
<ID>OUT</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>248</ID>
<type>GA_LED</type>
<position>25.5,-344</position>
<input>
<ID>N_in0</ID>121 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>249</ID>
<type>AA_LABEL</type>
<position>31,-297.5</position>
<gparam>LABEL_TEXT CARRY = AB </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>250</ID>
<type>AA_LABEL</type>
<position>40.5,-343</position>
<gparam>LABEL_TEXT CARRY = AB </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>252</ID>
<type>AA_LABEL</type>
<position>7.5,-356.5</position>
<gparam>LABEL_TEXT HALF SUBTRACTOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>253</ID>
<type>AA_AND2</type>
<position>5.5,-376.5</position>
<input>
<ID>IN_0</ID>128 </input>
<input>
<ID>IN_1</ID>127 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>254</ID>
<type>GA_LED</type>
<position>15,-376</position>
<input>
<ID>N_in0</ID>125 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>255</ID>
<type>AA_LABEL</type>
<position>28.5,-375</position>
<gparam>LABEL_TEXT B = AB </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>256</ID>
<type>AO_XNOR2</type>
<position>5,-367</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>127 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_TOGGLE</type>
<position>-14,-368</position>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>258</ID>
<type>AA_TOGGLE</type>
<position>-14.5,-373.5</position>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>259</ID>
<type>GA_LED</type>
<position>14.5,-367</position>
<input>
<ID>N_in0</ID>124 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>260</ID>
<type>AA_LABEL</type>
<position>-24,-367.5</position>
<gparam>LABEL_TEXT INPUT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>261</ID>
<type>AA_LABEL</type>
<position>-24,-373.5</position>
<gparam>LABEL_TEXT INPUT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>262</ID>
<type>AA_LABEL</type>
<position>17.5,-370</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>263</ID>
<type>AA_LABEL</type>
<position>32,-366.5</position>
<gparam>LABEL_TEXT D = AB + AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>264</ID>
<type>AA_LABEL</type>
<position>30,-363.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>265</ID>
<type>AA_LABEL</type>
<position>40,-363.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>267</ID>
<type>AE_SMALL_INVERTER</type>
<position>-7,-375.5</position>
<input>
<ID>IN_0</ID>126 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_LABEL</type>
<position>30,-372</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>269</ID>
<type>AA_LABEL</type>
<position>11,-386.5</position>
<gparam>LABEL_TEXT AOI IMPLIMENTATION</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>270</ID>
<type>AA_TOGGLE</type>
<position>-16,-398</position>
<output>
<ID>OUT_0</ID>139 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>271</ID>
<type>AA_TOGGLE</type>
<position>-4.5,-397.5</position>
<output>
<ID>OUT_0</ID>137 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>272</ID>
<type>AE_SMALL_INVERTER</type>
<position>-13,-402</position>
<input>
<ID>IN_0</ID>139 </input>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>273</ID>
<type>AE_SMALL_INVERTER</type>
<position>-1.5,-401</position>
<input>
<ID>IN_0</ID>137 </input>
<output>
<ID>OUT_0</ID>132 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>274</ID>
<type>AA_LABEL</type>
<position>-16,-394</position>
<gparam>LABEL_TEXT INPUT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>275</ID>
<type>AA_LABEL</type>
<position>-3.5,-394</position>
<gparam>LABEL_TEXT INPUT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>276</ID>
<type>AA_AND2</type>
<position>13,-406.5</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>137 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>277</ID>
<type>AA_AND2</type>
<position>12.5,-414.5</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>278</ID>
<type>AE_OR2</type>
<position>25,-409.5</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>134 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>GA_LED</type>
<position>33,-409.5</position>
<input>
<ID>N_in0</ID>135 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>280</ID>
<type>AA_AND2</type>
<position>12,-424.5</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>281</ID>
<type>GA_LED</type>
<position>24.5,-424.5</position>
<input>
<ID>N_in0</ID>136 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>287</ID>
<type>AA_LABEL</type>
<position>42.5,-421</position>
<gparam>LABEL_TEXT B = AB </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>288</ID>
<type>AA_LABEL</type>
<position>46,-412.5</position>
<gparam>LABEL_TEXT D = AB + AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>289</ID>
<type>AA_LABEL</type>
<position>44,-409.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>290</ID>
<type>AA_LABEL</type>
<position>54,-409.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>291</ID>
<type>AA_LABEL</type>
<position>44,-418</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>292</ID>
<type>AA_LABEL</type>
<position>12,-432</position>
<gparam>LABEL_TEXT NAND IMPLIMENTATION</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>AA_TOGGLE</type>
<position>-16,-439.5</position>
<output>
<ID>OUT_0</ID>149 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>294</ID>
<type>AA_TOGGLE</type>
<position>-2,-439.5</position>
<output>
<ID>OUT_0</ID>142 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>295</ID>
<type>BA_NAND2</type>
<position>-9.5,-444</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>149 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>296</ID>
<type>BA_NAND2</type>
<position>3.5,-444.5</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>142 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>297</ID>
<type>BA_NAND2</type>
<position>14.5,-452</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>141 </input>
<output>
<ID>OUT</ID>144 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>298</ID>
<type>BA_NAND2</type>
<position>15,-460.5</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>299</ID>
<type>BA_NAND2</type>
<position>26.5,-456</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>300</ID>
<type>GA_LED</type>
<position>34.5,-456</position>
<input>
<ID>N_in0</ID>146 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>305</ID>
<type>BA_NAND2</type>
<position>15.5,-471</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>142 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>306</ID>
<type>BA_NAND2</type>
<position>30,-471</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>147 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>307</ID>
<type>GA_LED</type>
<position>37,-471</position>
<input>
<ID>N_in0</ID>148 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>309</ID>
<type>AA_LABEL</type>
<position>46.5,-465.5</position>
<gparam>LABEL_TEXT B = AB </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>310</ID>
<type>AA_LABEL</type>
<position>50,-457</position>
<gparam>LABEL_TEXT D = AB + AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>311</ID>
<type>AA_LABEL</type>
<position>48,-454</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>312</ID>
<type>AA_LABEL</type>
<position>58,-454</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>313</ID>
<type>AA_LABEL</type>
<position>48,-462.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>314</ID>
<type>AA_LABEL</type>
<position>-14.5,-436</position>
<gparam>LABEL_TEXT INPUT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>315</ID>
<type>AA_LABEL</type>
<position>-2,-436</position>
<gparam>LABEL_TEXT INPUT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,43,-29,43</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-41 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>-41,43,-41,45</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>43 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,41,-29,41</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-41 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-41,39,-41,41</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>41 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-23,42,-21,42</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>-21 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>-21,41.5,-21,42</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<intersection>42 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-35,27.5,-29.5,27.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-35 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-35,27.5,-35,29.5</points>
<intersection>27.5 1</intersection>
<intersection>29.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-41,29.5,-35,29.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-35 5</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,24,-35.5,25.5</points>
<intersection>24 2</intersection>
<intersection>25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35.5,25.5,-29.5,25.5</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>-35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-41,24,-35.5,24</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>-35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-23.5,26.5,-20.5,26.5</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<connection>
<GID>27</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,12.5,-35.5,13.5</points>
<intersection>12.5 1</intersection>
<intersection>13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35.5,12.5,-29.5,12.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>-35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-42,13.5,-35.5,13.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>-35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,8.5,-35.5,10.5</points>
<intersection>8.5 2</intersection>
<intersection>10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35.5,10.5,-29.5,10.5</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>-35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-42,8.5,-35.5,8.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-23.5,11.5,-21,11.5</points>
<connection>
<GID>38</GID>
<name>N_in0</name></connection>
<connection>
<GID>36</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-5,-36,-3</points>
<intersection>-5 1</intersection>
<intersection>-3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-5,-29.5,-5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-42,-3,-36,-3</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-9,-36,-7</points>
<intersection>-9 2</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-7,-29.5,-7</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-42,-9,-36,-9</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-23.5,-6,-22,-6</points>
<connection>
<GID>51</GID>
<name>N_in0</name></connection>
<connection>
<GID>49</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,44.5,27.5,45.5</points>
<intersection>44.5 1</intersection>
<intersection>45.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,44.5,35.5,44.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,45.5,27.5,45.5</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,40.5,27.5,42.5</points>
<intersection>40.5 2</intersection>
<intersection>42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,42.5,35.5,42.5</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,40.5,27.5,40.5</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41.5,43.5,46.5,43.5</points>
<connection>
<GID>61</GID>
<name>N_in0</name></connection>
<connection>
<GID>63</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10,-32,-4,-32</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>-4 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-4,-33,-4,-31</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>-32 1</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2,-32,6,-32</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<connection>
<GID>76</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-40.5,-7,-40</points>
<intersection>-40.5 1</intersection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,-40.5,-4,-40.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>-7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-10,-40,-7,-40</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-44,-7,-42.5</points>
<intersection>-44 2</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,-42.5,-4,-42.5</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>-7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-10,-44,-7,-44</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2,-41.5,7,-41.5</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>6 4</intersection>
<intersection>7 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>6,-42.5,6,-41.5</points>
<intersection>-42.5 5</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>6,-42.5,7,-42.5</points>
<connection>
<GID>84</GID>
<name>IN_1</name></connection>
<intersection>6 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>7,-41.5,7,-40.5</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>-41.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-41.5,16.5,-41.5</points>
<connection>
<GID>85</GID>
<name>N_in0</name></connection>
<connection>
<GID>84</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10,-51.5,-4.5,-51.5</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<intersection>-4.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-4.5,-52.5,-4.5,-50.5</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>-51.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10,-59,-4.5,-59</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>-4.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-4.5,-60,-4.5,-58</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>-59 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-54,3.5,-51.5</points>
<intersection>-54 1</intersection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,-54,6,-54</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1.5,-51.5,3.5,-51.5</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-59,3.5,-56</points>
<intersection>-59 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,-56,6,-56</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1.5,-59,3.5,-59</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,-55,16,-55</points>
<connection>
<GID>92</GID>
<name>N_in0</name></connection>
<connection>
<GID>91</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-4,-69,-4,-67</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>-68 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-10,-68,-4,-68</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<intersection>-4 3</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-4,-77.5,-4,-75.5</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>-76.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-10,-76.5,-4,-76.5</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<intersection>-4 3</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>16,-72.5,16,-70.5</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>-71.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>12.5,-71.5,16,-71.5</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<intersection>16 3</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-71.5,26.5,-71.5</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<connection>
<GID>100</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-70.5,4,-68</points>
<intersection>-70.5 1</intersection>
<intersection>-68 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-70.5,6.5,-70.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2,-68,4,-68</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<intersection>4 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-76.5,4,-72.5</points>
<intersection>-76.5 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-72.5,6.5,-72.5</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2,-76.5,4,-76.5</points>
<connection>
<GID>95</GID>
<name>OUT</name></connection>
<intersection>4 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10,-85,4.5,-85</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-10 6</intersection>
<intersection>-7 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-7,-88.5,-7,-85</points>
<intersection>-88.5 5</intersection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-7,-88.5,-5,-88.5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>-7 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-10,-85.5,-10,-85</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>-85 1</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10,-93.5,5,-93.5</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>-7 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-7,-93.5,-7,-90.5</points>
<intersection>-93.5 1</intersection>
<intersection>-90.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-7,-90.5,-5,-90.5</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>-7 4</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-91.5,2.5,-87</points>
<intersection>-91.5 3</intersection>
<intersection>-89.5 2</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,-87,4.5,-87</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1,-89.5,2.5,-89.5</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>2.5,-91.5,5,-91.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-88,12.5,-86</points>
<intersection>-88 1</intersection>
<intersection>-86 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12.5,-88,14.5,-88</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10.5,-86,12.5,-86</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-92.5,13,-90</points>
<intersection>-92.5 2</intersection>
<intersection>-90 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-90,14.5,-90</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-92.5,13,-92.5</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>13 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-89,25.5,-89</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<connection>
<GID>116</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10,-101.5,4.5,-101.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>-10 6</intersection>
<intersection>-7 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-7,-105,-7,-101.5</points>
<intersection>-105 5</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-7,-105,-5,-105</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>-7 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-10,-102,-10,-101.5</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>-101.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10,-110,5,-110</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>-7 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-7,-110,-7,-107</points>
<intersection>-110 1</intersection>
<intersection>-107 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-7,-107,-5,-107</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>-7 4</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-108,2.5,-103.5</points>
<intersection>-108 3</intersection>
<intersection>-106 2</intersection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,-103.5,4.5,-103.5</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1,-106,2.5,-106</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>2.5,-108,5,-108</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-104.5,12.5,-102.5</points>
<intersection>-104.5 1</intersection>
<intersection>-102.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12.5,-104.5,14.5,-104.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10.5,-102.5,12.5,-102.5</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-109,13,-106.5</points>
<intersection>-109 2</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-106.5,14.5,-106.5</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-109,13,-109</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<intersection>13 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-106.5,21.5,-104.5</points>
<intersection>-106.5 3</intersection>
<intersection>-105.5 2</intersection>
<intersection>-104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-104.5,23,-104.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20.5,-105.5,21.5,-105.5</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>21.5,-106.5,23,-106.5</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-105.5,32.5,-105.5</points>
<connection>
<GID>124</GID>
<name>N_in0</name></connection>
<connection>
<GID>125</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-10.5,-137.5,-5.5,-137.5</points>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<intersection>-5.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-5.5,-138.5,-5.5,-136.5</points>
<intersection>-138.5 5</intersection>
<intersection>-137.5 1</intersection>
<intersection>-136.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-5.5,-136.5,-4.5,-136.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-5.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-5.5,-138.5,-4.5,-138.5</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>-5.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>1.5,-137.5,2.5,-137.5</points>
<connection>
<GID>133</GID>
<name>N_in0</name></connection>
<connection>
<GID>130</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-146.5,-7.5,-145.5</points>
<intersection>-146.5 1</intersection>
<intersection>-145.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-146.5,-5,-146.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-10.5,-145.5,-7.5,-145.5</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-150,-7.5,-148.5</points>
<intersection>-150 2</intersection>
<intersection>-148.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-148.5,-5,-148.5</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-10.5,-150,-7.5,-150</points>
<connection>
<GID>137</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>4,-148.5,4,-146.5</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>-147.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>1,-147.5,4,-147.5</points>
<connection>
<GID>135</GID>
<name>OUT</name></connection>
<intersection>4 3</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-147.5,12,-147.5</points>
<connection>
<GID>141</GID>
<name>N_in0</name></connection>
<connection>
<GID>140</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11,-159,-6,-159</points>
<connection>
<GID>145</GID>
<name>OUT_0</name></connection>
<intersection>-6 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-6,-160,-6,-158</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>-159 1</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11,-166,-6,-166</points>
<connection>
<GID>147</GID>
<name>OUT_0</name></connection>
<intersection>-6 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-6,-167,-6,-165</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>-166 1</intersection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9.5,-162.5,12.5,-162.5</points>
<connection>
<GID>149</GID>
<name>N_in0</name></connection>
<intersection>9.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>9.5,-162.5,9.5,-162.5</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<intersection>-162.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-161.5,2,-159</points>
<intersection>-161.5 1</intersection>
<intersection>-159 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-161.5,3.5,-161.5</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0,-159,2,-159</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-166,2,-163.5</points>
<intersection>-166 2</intersection>
<intersection>-163.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-163.5,3.5,-163.5</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0,-166,2,-166</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11,-176.5,-6,-176.5</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>-6 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-6,-177.5,-6,-175.5</points>
<connection>
<GID>151</GID>
<name>IN_1</name></connection>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>-176.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11,-183.5,-6,-183.5</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<intersection>-6 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-6,-184.5,-6,-182.5</points>
<connection>
<GID>153</GID>
<name>IN_1</name></connection>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>-183.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-179,2,-176.5</points>
<intersection>-179 1</intersection>
<intersection>-176.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-179,3.5,-179</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0,-176.5,2,-176.5</points>
<connection>
<GID>151</GID>
<name>OUT</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-183.5,2,-181</points>
<intersection>-183.5 2</intersection>
<intersection>-181 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-181,3.5,-181</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0,-183.5,2,-183.5</points>
<connection>
<GID>153</GID>
<name>OUT</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-181,11,-179</points>
<intersection>-181 3</intersection>
<intersection>-180 2</intersection>
<intersection>-179 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-179,12.5,-179</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-180,11,-180</points>
<connection>
<GID>155</GID>
<name>OUT</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>11,-181,12.5,-181</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,-180,20.5,-180</points>
<connection>
<GID>157</GID>
<name>N_in0</name></connection>
<connection>
<GID>156</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-197.5,-9.5,-192</points>
<intersection>-197.5 5</intersection>
<intersection>-194.5 2</intersection>
<intersection>-192 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9.5,-192,1,-192</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-12.5,-194.5,-9.5,-194.5</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-9.5,-197.5,-7,-197.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>-9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-205,-9.5,-199.5</points>
<intersection>-205 4</intersection>
<intersection>-203 2</intersection>
<intersection>-199.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9.5,-199.5,-7,-199.5</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-12.5,-203,-9.5,-203</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-9.5,-205,1,-205</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<intersection>-9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,-203,0,-194</points>
<intersection>-203 3</intersection>
<intersection>-198.5 2</intersection>
<intersection>-194 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-194,1,-194</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>0 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1,-198.5,0,-198.5</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<intersection>0 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>0,-203,1,-203</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>0 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-197,8.5,-193</points>
<intersection>-197 1</intersection>
<intersection>-193 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-197,10.5,-197</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-193,8.5,-193</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-204,8.5,-199</points>
<intersection>-204 2</intersection>
<intersection>-199 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-199,10.5,-199</points>
<connection>
<GID>165</GID>
<name>IN_1</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-204,8.5,-204</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>18.5,-199,18.5,-197</points>
<intersection>-199 5</intersection>
<intersection>-198 6</intersection>
<intersection>-197 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>18.5,-197,19.5,-197</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>18.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>18.5,-199,19.5,-199</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<intersection>18.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>16.5,-198,18.5,-198</points>
<connection>
<GID>165</GID>
<name>OUT</name></connection>
<intersection>18.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>25.5,-198,26.5,-198</points>
<connection>
<GID>167</GID>
<name>N_in0</name></connection>
<connection>
<GID>166</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-218.5,-9.5,-213</points>
<intersection>-218.5 5</intersection>
<intersection>-215 2</intersection>
<intersection>-213 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9.5,-213,1,-213</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-13.5,-215,-9.5,-215</points>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-9.5,-218.5,-7,-218.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>-9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-226,-9.5,-220.5</points>
<intersection>-226 4</intersection>
<intersection>-223.5 2</intersection>
<intersection>-220.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9.5,-220.5,-7,-220.5</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-14.5,-223.5,-9.5,-223.5</points>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-9.5,-226,1,-226</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>-9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,-224,0,-215</points>
<intersection>-224 3</intersection>
<intersection>-219.5 2</intersection>
<intersection>-215 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-215,1,-215</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>0 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1,-219.5,0,-219.5</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<intersection>0 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>0,-224,1,-224</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>0 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-218,8.5,-214</points>
<intersection>-218 1</intersection>
<intersection>-214 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-218,10.5,-218</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-214,8.5,-214</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-225,8.5,-220</points>
<intersection>-225 2</intersection>
<intersection>-220 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-220,10.5,-220</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-225,8.5,-225</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-219,20.5,-219</points>
<connection>
<GID>176</GID>
<name>N_in0</name></connection>
<connection>
<GID>174</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-9.5,-249.5,-7,-249.5</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>-9.5 4</intersection>
<intersection>-7.5 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-9.5,-249.5,-9.5,-248</points>
<intersection>-249.5 1</intersection>
<intersection>-248 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-12.5,-248,-9.5,-248</points>
<connection>
<GID>182</GID>
<name>OUT_0</name></connection>
<intersection>-9.5 4</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-7.5,-256.5,-7.5,-249.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>-249.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-258.5,-9.5,-251.5</points>
<intersection>-258.5 3</intersection>
<intersection>-253.5 2</intersection>
<intersection>-251.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9.5,-251.5,-7,-251.5</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-12.5,-253.5,-9.5,-253.5</points>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-9.5,-258.5,-7.5,-258.5</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>-9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-250.5,3,-250.5</points>
<connection>
<GID>184</GID>
<name>N_in0</name></connection>
<connection>
<GID>181</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-257.5,2.5,-257.5</points>
<connection>
<GID>200</GID>
<name>N_in0</name></connection>
<connection>
<GID>198</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21.5,-279,-21.5,-275.5</points>
<intersection>-279 1</intersection>
<intersection>-275.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21.5,-279,-1.5,-279</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-22.5,-275.5,-21.5,-275.5</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<intersection>-21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-297,-16,-273</points>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection>
<intersection>-297 5</intersection>
<intersection>-281 1</intersection>
<intersection>-274.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-281,-1.5,-281</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-16,-274.5,-15,-274.5</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-16,-297,-2.5,-297</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27.5,-299,-27.5,-273</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>-299 5</intersection>
<intersection>-286.5 1</intersection>
<intersection>-275.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27.5,-286.5,-1.5,-286.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>-27.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-27.5,-275.5,-26.5,-275.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>-27.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-27.5,-299,-2.5,-299</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>-27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-288.5,-10,-274.5</points>
<intersection>-288.5 1</intersection>
<intersection>-274.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10,-288.5,-1.5,-288.5</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-11,-274.5,-10,-274.5</points>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-282,7.5,-280</points>
<intersection>-282 1</intersection>
<intersection>-280 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,-282,10.5,-282</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-280,7.5,-280</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-287.5,7.5,-284</points>
<intersection>-287.5 1</intersection>
<intersection>-284 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4.5,-287.5,7.5,-287.5</points>
<connection>
<GID>213</GID>
<name>OUT</name></connection>
<intersection>7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-284,10.5,-284</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-283,20.5,-283</points>
<connection>
<GID>217</GID>
<name>N_in0</name></connection>
<connection>
<GID>215</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-298,12,-298</points>
<connection>
<GID>221</GID>
<name>N_in0</name></connection>
<connection>
<GID>219</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27.5,-343,-27.5,-314.5</points>
<connection>
<GID>229</GID>
<name>OUT_0</name></connection>
<intersection>-343 5</intersection>
<intersection>-324 1</intersection>
<intersection>-317 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27.5,-324,0,-324</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>-27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27.5,-317,-24,-317</points>
<intersection>-27.5 0</intersection>
<intersection>-24 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-24,-318,-24,-316</points>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>-317 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-27.5,-343,1,-343</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>-27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-326,-4.5,-317.5</points>
<intersection>-326 1</intersection>
<intersection>-317.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-326,0,-326</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-5,-317.5,-4.5,-317.5</points>
<connection>
<GID>235</GID>
<name>OUT</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-345,-13.5,-314.5</points>
<connection>
<GID>231</GID>
<name>OUT_0</name></connection>
<intersection>-345 5</intersection>
<intersection>-332.5 1</intersection>
<intersection>-317 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13.5,-332.5,0.5,-332.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>-13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-13.5,-317,-11,-317</points>
<intersection>-13.5 0</intersection>
<intersection>-11 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-11,-318.5,-11,-316.5</points>
<connection>
<GID>235</GID>
<name>IN_1</name></connection>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>-317 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-13.5,-345,1,-345</points>
<connection>
<GID>245</GID>
<name>IN_1</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17.5,-334.5,-17.5,-317</points>
<intersection>-334.5 1</intersection>
<intersection>-317 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17.5,-334.5,0.5,-334.5</points>
<connection>
<GID>237</GID>
<name>IN_1</name></connection>
<intersection>-17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-18,-317,-17.5,-317</points>
<connection>
<GID>233</GID>
<name>OUT</name></connection>
<intersection>-17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-328,9,-325</points>
<intersection>-328 1</intersection>
<intersection>-325 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-328,12,-328</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-325,9,-325</points>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-333.5,9,-330</points>
<intersection>-333.5 2</intersection>
<intersection>-330 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-330,12,-330</points>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-333.5,9,-333.5</points>
<connection>
<GID>237</GID>
<name>OUT</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-329,22,-329</points>
<connection>
<GID>239</GID>
<name>N_in0</name></connection>
<connection>
<GID>238</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-344,14.5,-344</points>
<connection>
<GID>245</GID>
<name>OUT</name></connection>
<intersection>14.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>14.5,-345,14.5,-343</points>
<intersection>-345 6</intersection>
<intersection>-344 1</intersection>
<intersection>-343 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>14.5,-343,15.5,-343</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>14.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>14.5,-345,15.5,-345</points>
<connection>
<GID>247</GID>
<name>IN_1</name></connection>
<intersection>14.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-344,24.5,-344</points>
<connection>
<GID>248</GID>
<name>N_in0</name></connection>
<connection>
<GID>247</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8,-367,13.5,-367</points>
<connection>
<GID>256</GID>
<name>OUT</name></connection>
<connection>
<GID>259</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-376.5,14,-376.5</points>
<connection>
<GID>253</GID>
<name>OUT</name></connection>
<intersection>14 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>14,-376.5,14,-376</points>
<connection>
<GID>254</GID>
<name>N_in0</name></connection>
<intersection>-376.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-368,-5,-366</points>
<intersection>-368 2</intersection>
<intersection>-366 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-366,2,-366</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-12,-368,-5,-368</points>
<connection>
<GID>257</GID>
<name>OUT_0</name></connection>
<intersection>-9 3</intersection>
<intersection>-5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-9,-375.5,-9,-368</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>-368 2</intersection></vsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10.5,-377.5,-10.5,-370.5</points>
<intersection>-377.5 3</intersection>
<intersection>-373.5 2</intersection>
<intersection>-370.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10.5,-370.5,2,-370.5</points>
<intersection>-10.5 0</intersection>
<intersection>2 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-12.5,-373.5,-10.5,-373.5</points>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<intersection>-10.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-10.5,-377.5,2.5,-377.5</points>
<connection>
<GID>253</GID>
<name>IN_1</name></connection>
<intersection>-10.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>2,-370.5,2,-368</points>
<connection>
<GID>256</GID>
<name>IN_1</name></connection>
<intersection>-370.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5,-375.5,2.5,-375.5</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-425.5,-10,-402</points>
<intersection>-425.5 4</intersection>
<intersection>-405.5 1</intersection>
<intersection>-402 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10,-405.5,10,-405.5</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-11,-402,-10,-402</points>
<connection>
<GID>272</GID>
<name>OUT_0</name></connection>
<intersection>-10 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-10,-425.5,9,-425.5</points>
<connection>
<GID>280</GID>
<name>IN_1</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1.5,-415.5,1.5,-401</points>
<intersection>-415.5 1</intersection>
<intersection>-401 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1.5,-415.5,9.5,-415.5</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0.5,-401,1.5,-401</points>
<connection>
<GID>273</GID>
<name>OUT_0</name></connection>
<intersection>1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-408.5,19,-406.5</points>
<intersection>-408.5 1</intersection>
<intersection>-406.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-408.5,22,-408.5</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-406.5,19,-406.5</points>
<connection>
<GID>276</GID>
<name>OUT</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-414.5,19,-410.5</points>
<intersection>-414.5 1</intersection>
<intersection>-410.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,-414.5,19,-414.5</points>
<connection>
<GID>277</GID>
<name>OUT</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,-410.5,22,-410.5</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-409.5,32,-409.5</points>
<connection>
<GID>279</GID>
<name>N_in0</name></connection>
<connection>
<GID>278</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-424.5,23.5,-424.5</points>
<connection>
<GID>281</GID>
<name>N_in0</name></connection>
<connection>
<GID>280</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-423.5,-4.5,-399.5</points>
<connection>
<GID>271</GID>
<name>OUT_0</name></connection>
<intersection>-423.5 1</intersection>
<intersection>-407.5 3</intersection>
<intersection>-401 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-423.5,9,-423.5</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4.5,-401,-3.5,-401</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-407.5,10,-407.5</points>
<connection>
<GID>276</GID>
<name>IN_1</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-413.5,-16,-400</points>
<connection>
<GID>270</GID>
<name>OUT_0</name></connection>
<intersection>-413.5 1</intersection>
<intersection>-402 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-413.5,9.5,-413.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-16,-402,-15,-402</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-453,7,-444.5</points>
<intersection>-453 1</intersection>
<intersection>-444.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7,-453,11.5,-453</points>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-444.5,7,-444.5</points>
<connection>
<GID>296</GID>
<name>OUT</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-472,-2,-441.5</points>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection>
<intersection>-472 5</intersection>
<intersection>-459.5 1</intersection>
<intersection>-444 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2,-459.5,12,-459.5</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,-444,0.5,-444</points>
<intersection>-2 0</intersection>
<intersection>0.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>0.5,-445.5,0.5,-443.5</points>
<connection>
<GID>296</GID>
<name>IN_1</name></connection>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>-444 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-2,-472,12.5,-472</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-455,20.5,-452</points>
<intersection>-455 1</intersection>
<intersection>-452 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-455,23.5,-455</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-452,20.5,-452</points>
<connection>
<GID>297</GID>
<name>OUT</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-460.5,20.5,-457</points>
<intersection>-460.5 2</intersection>
<intersection>-457 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-457,23.5,-457</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-460.5,20.5,-460.5</points>
<connection>
<GID>298</GID>
<name>OUT</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-456,33.5,-456</points>
<connection>
<GID>300</GID>
<name>N_in0</name></connection>
<connection>
<GID>299</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,-471,26,-471</points>
<connection>
<GID>305</GID>
<name>OUT</name></connection>
<intersection>26 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>26,-472,26,-470</points>
<intersection>-472 6</intersection>
<intersection>-471 1</intersection>
<intersection>-470 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>26,-470,27,-470</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>26 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>26,-472,27,-472</points>
<connection>
<GID>306</GID>
<name>IN_1</name></connection>
<intersection>26 4</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33,-471,36,-471</points>
<connection>
<GID>307</GID>
<name>N_in0</name></connection>
<connection>
<GID>306</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-451,-16,-441.5</points>
<connection>
<GID>293</GID>
<name>OUT_0</name></connection>
<intersection>-451 1</intersection>
<intersection>-444 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-451,11.5,-451</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-16,-444,-12.5,-444</points>
<intersection>-16 0</intersection>
<intersection>-12.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-12.5,-445,-12.5,-443</points>
<connection>
<GID>295</GID>
<name>IN_1</name></connection>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>-444 2</intersection></vsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-470,-6,-444</points>
<intersection>-470 4</intersection>
<intersection>-461.5 1</intersection>
<intersection>-444 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-461.5,12,-461.5</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<intersection>-6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-6.5,-444,-6,-444</points>
<connection>
<GID>295</GID>
<name>OUT</name></connection>
<intersection>-6 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-6,-470,12.5,-470</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 9></circuit>