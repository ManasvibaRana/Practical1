<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-187.67,-6.23354,311.32,-252.875</PageViewport>
<gate>
<ID>2</ID>
<type>BA_NAND2</type>
<position>33.5,-16</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>17.5,-8</position>
<gparam>LABEL_TEXT SR latch NAND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>BA_NAND2</type>
<position>33.5,-25</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>43,-16</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>43,-25</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>19.5,-15</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>20,-26</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>17,-14.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>17.5,-25.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>46,-15.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>46,-25</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>46,-22</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>93.5,-16</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>93.5,-25</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>71,-14.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>70.5,-26</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>68,-25.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>67.5,-15</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>96.5,-15.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>96.5,-25</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>96.5,-22</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>73,-7</position>
<gparam>LABEL_TEXT SR latch NOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>BE_NOR2</type>
<position>83.5,-15.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>BE_NOR2</type>
<position>83.5,-26</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>16.5,-34.5</position>
<gparam>LABEL_TEXT SR Flip Flop</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>BA_NAND2</type>
<position>35,-47.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>BA_NAND2</type>
<position>35,-56.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>GA_LED</type>
<position>44.5,-47.5</position>
<input>
<ID>N_in0</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>GA_LED</type>
<position>44.5,-56.5</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_TOGGLE</type>
<position>9,-46</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>8.5,-57</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>5.5,-46</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>5,-56.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>47.5,-47</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>47.5,-56.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>47.5,-53.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>BA_NAND2</type>
<position>20,-46.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>BA_NAND2</type>
<position>21,-57.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>BB_CLOCK</type>
<position>12.5,-51</position>
<output>
<ID>CLK</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>68</ID>
<type>BA_NAND2</type>
<position>98.5,-47.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>BA_NAND2</type>
<position>98.5,-56.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>GA_LED</type>
<position>108,-47.5</position>
<input>
<ID>N_in0</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>GA_LED</type>
<position>108,-56.5</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>70.5,-42.5</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>70.5,-40</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>111,-47</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>111,-56.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>111,-54</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>BA_NAND2</type>
<position>83.5,-46.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>BA_NAND2</type>
<position>84.5,-57.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>BB_CLOCK</type>
<position>76,-51</position>
<output>
<ID>CLK</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_LABEL</type>
<position>74.5,-35.5</position>
<gparam>LABEL_TEXT D Flip Flop</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AE_SMALL_INVERTER</type>
<position>70.5,-50</position>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>86</ID>
<type>AE_DFF_LOW</type>
<position>86,-70</position>
<input>
<ID>IN_0</ID>37 </input>
<output>
<ID>OUTINV_0</ID>39 </output>
<output>
<ID>OUT_0</ID>38 </output>
<input>
<ID>clock</ID>36 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>88</ID>
<type>BB_CLOCK</type>
<position>78,-71</position>
<output>
<ID>CLK</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_TOGGLE</type>
<position>77.5,-66.5</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>92</ID>
<type>GA_LED</type>
<position>93,-68</position>
<input>
<ID>N_in0</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>GA_LED</type>
<position>93.5,-71</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>21.5,-83.5</position>
<gparam>LABEL_TEXT JK Flip Flop</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>BE_JKFF_LOW</type>
<position>41,-95</position>
<input>
<ID>J</ID>48 </input>
<input>
<ID>K</ID>49 </input>
<output>
<ID>Q</ID>50 </output>
<input>
<ID>clock</ID>47 </input>
<output>
<ID>nQ</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>113</ID>
<type>BB_CLOCK</type>
<position>31,-95</position>
<output>
<ID>CLK</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_TOGGLE</type>
<position>30,-90.5</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_TOGGLE</type>
<position>31,-99</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>119</ID>
<type>GA_LED</type>
<position>48.5,-93</position>
<input>
<ID>N_in0</ID>50 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>GA_LED</type>
<position>48.5,-97</position>
<input>
<ID>N_in0</ID>51 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>51.5,-97</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>51.5,-94.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_LABEL</type>
<position>51.5,-92.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>AA_LABEL</type>
<position>27.5,-90</position>
<gparam>LABEL_TEXT J</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>27.5,-99</position>
<gparam>LABEL_TEXT K</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>AA_LABEL</type>
<position>81,-80.5</position>
<gparam>LABEL_TEXT T Flip Flop</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>BE_JKFF_LOW</type>
<position>91.5,-96</position>
<input>
<ID>J</ID>67 </input>
<input>
<ID>K</ID>67 </input>
<output>
<ID>Q</ID>65 </output>
<input>
<ID>clock</ID>62 </input>
<output>
<ID>nQ</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>153</ID>
<type>BB_CLOCK</type>
<position>81.5,-96</position>
<output>
<ID>CLK</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>154</ID>
<type>AA_TOGGLE</type>
<position>76,-88</position>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>156</ID>
<type>GA_LED</type>
<position>99,-94</position>
<input>
<ID>N_in0</ID>65 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>GA_LED</type>
<position>99,-98</position>
<input>
<ID>N_in0</ID>66 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>AA_LABEL</type>
<position>102,-98</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>AA_LABEL</type>
<position>102,-95.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>AA_LABEL</type>
<position>102,-93.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>76,-85.5</position>
<gparam>LABEL_TEXT T</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>AA_LABEL</type>
<position>19,-106</position>
<gparam>LABEL_TEXT D TO SR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>AE_DFF_LOW</type>
<position>35.5,-122.5</position>
<input>
<ID>IN_0</ID>76 </input>
<output>
<ID>OUTINV_0</ID>69 </output>
<output>
<ID>OUT_0</ID>73 </output>
<input>
<ID>clock</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>167</ID>
<type>GA_LED</type>
<position>52,-121</position>
<input>
<ID>N_in0</ID>73 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>GA_LED</type>
<position>51,-125.5</position>
<input>
<ID>N_in0</ID>69 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>AA_TOGGLE</type>
<position>18.5,-113</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>173</ID>
<type>BB_CLOCK</type>
<position>26,-136.5</position>
<output>
<ID>CLK</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_TOGGLE</type>
<position>14.5,-113</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>177</ID>
<type>AE_SMALL_INVERTER</type>
<position>18.5,-118</position>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_AND2</type>
<position>19.5,-124</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>181</ID>
<type>AE_OR2</type>
<position>15.5,-130.5</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_LABEL</type>
<position>54.5,-125.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_LABEL</type>
<position>54.5,-123</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>54.5,-121</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>AA_LABEL</type>
<position>14.5,-110</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>18.5,-110</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>BA_NAND2</type>
<position>96.5,-142</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>BA_NAND2</type>
<position>96.5,-151</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>GA_LED</type>
<position>106,-142</position>
<input>
<ID>N_in0</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>GA_LED</type>
<position>106,-151</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>193</ID>
<type>AA_LABEL</type>
<position>109,-141.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>194</ID>
<type>AA_LABEL</type>
<position>109,-151</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>195</ID>
<type>AA_LABEL</type>
<position>109,-148.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>196</ID>
<type>BA_NAND2</type>
<position>81.5,-141</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>197</ID>
<type>BA_NAND2</type>
<position>82.5,-152</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>198</ID>
<type>BB_CLOCK</type>
<position>74,-145.5</position>
<output>
<ID>CLK</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>199</ID>
<type>AE_SMALL_INVERTER</type>
<position>68.5,-144.5</position>
<input>
<ID>IN_0</ID>82 </input>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_TOGGLE</type>
<position>52.5,-134</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_TOGGLE</type>
<position>56.5,-134</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>202</ID>
<type>AE_SMALL_INVERTER</type>
<position>57,-139</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>203</ID>
<type>AA_AND2</type>
<position>58,-145</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>204</ID>
<type>AE_OR2</type>
<position>54,-151.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_LABEL</type>
<position>52.5,-131</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>206</ID>
<type>AA_LABEL</type>
<position>56.5,-131</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>207</ID>
<type>AA_LABEL</type>
<position>14.5,-160</position>
<gparam>LABEL_TEXT D TO JK</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AE_DFF_LOW</type>
<position>36,-176</position>
<input>
<ID>IN_0</ID>97 </input>
<output>
<ID>OUTINV_0</ID>89 </output>
<output>
<ID>OUT_0</ID>88 </output>
<input>
<ID>clock</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_TOGGLE</type>
<position>11,-172.5</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>213</ID>
<type>AA_TOGGLE</type>
<position>11,-179.5</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>215</ID>
<type>BB_CLOCK</type>
<position>25.5,-190</position>
<output>
<ID>CLK</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>217</ID>
<type>GA_LED</type>
<position>47,-174</position>
<input>
<ID>N_in0</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>GA_LED</type>
<position>47,-177.5</position>
<input>
<ID>N_in0</ID>89 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>221</ID>
<type>AA_AND2</type>
<position>18.5,-171.5</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>92 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>223</ID>
<type>AE_SMALL_INVERTER</type>
<position>16,-179.5</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>225</ID>
<type>AA_AND2</type>
<position>21.5,-180.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>AE_OR2</type>
<position>27.5,-174.5</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>AA_LABEL</type>
<position>50,-173.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>231</ID>
<type>AA_LABEL</type>
<position>50,-177.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>AA_LABEL</type>
<position>50,-175</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>233</ID>
<type>AA_LABEL</type>
<position>8,-172</position>
<gparam>LABEL_TEXT J</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>237</ID>
<type>AA_LABEL</type>
<position>8.5,-179</position>
<gparam>LABEL_TEXT K</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>238</ID>
<type>AA_LABEL</type>
<position>76.5,-160</position>
<gparam>LABEL_TEXT D TO T</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>240</ID>
<type>AE_DFF_LOW</type>
<position>86,-176.5</position>
<input>
<ID>IN_0</ID>102 </input>
<output>
<ID>OUTINV_0</ID>99 </output>
<output>
<ID>OUT_0</ID>98 </output>
<input>
<ID>clock</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>241</ID>
<type>GA_LED</type>
<position>93.5,-174.5</position>
<input>
<ID>N_in0</ID>98 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>GA_LED</type>
<position>93.5,-178</position>
<input>
<ID>N_in0</ID>99 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>243</ID>
<type>AA_LABEL</type>
<position>96.5,-174</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>244</ID>
<type>AA_LABEL</type>
<position>96.5,-178</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>AA_LABEL</type>
<position>96.5,-175.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>246</ID>
<type>BB_CLOCK</type>
<position>77,-183</position>
<output>
<ID>CLK</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>247</ID>
<type>AA_TOGGLE</type>
<position>66.5,-173</position>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>249</ID>
<type>AI_XOR2</type>
<position>75,-172.5</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_LABEL</type>
<position>64,-172.5</position>
<gparam>LABEL_TEXT T</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>251</ID>
<type>AA_LABEL</type>
<position>16,-201</position>
<gparam>LABEL_TEXT JK TO SR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>253</ID>
<type>BE_JKFF_LOW</type>
<position>29.5,-215.5</position>
<input>
<ID>J</ID>103 </input>
<input>
<ID>K</ID>104 </input>
<output>
<ID>Q</ID>106 </output>
<input>
<ID>clock</ID>105 </input>
<output>
<ID>nQ</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_TOGGLE</type>
<position>15.5,-212</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_TOGGLE</type>
<position>15.5,-220</position>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>259</ID>
<type>BB_CLOCK</type>
<position>19,-215.5</position>
<output>
<ID>CLK</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>261</ID>
<type>GA_LED</type>
<position>36.5,-213</position>
<input>
<ID>N_in0</ID>106 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>263</ID>
<type>GA_LED</type>
<position>36.5,-217.5</position>
<input>
<ID>N_in0</ID>107 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>264</ID>
<type>AA_LABEL</type>
<position>53.5,-200.5</position>
<gparam>LABEL_TEXT JK TO D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>266</ID>
<type>AA_LABEL</type>
<position>13,-211.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>267</ID>
<type>AA_LABEL</type>
<position>12.5,-219.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>268</ID>
<type>AA_LABEL</type>
<position>39.5,-213</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>269</ID>
<type>AA_LABEL</type>
<position>39.5,-217</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>270</ID>
<type>AA_LABEL</type>
<position>39.5,-214.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>286</ID>
<type>BE_JKFF_LOW</type>
<position>67,-214</position>
<input>
<ID>J</ID>114 </input>
<input>
<ID>K</ID>115 </input>
<output>
<ID>Q</ID>116 </output>
<input>
<ID>clock</ID>113 </input>
<output>
<ID>nQ</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>287</ID>
<type>BB_CLOCK</type>
<position>54.5,-214</position>
<output>
<ID>CLK</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>288</ID>
<type>AA_TOGGLE</type>
<position>49,-207</position>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>289</ID>
<type>AE_SMALL_INVERTER</type>
<position>49,-214.5</position>
<input>
<ID>IN_0</ID>114 </input>
<output>
<ID>OUT_0</ID>115 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>290</ID>
<type>GA_LED</type>
<position>74.5,-212</position>
<input>
<ID>N_in0</ID>116 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>291</ID>
<type>GA_LED</type>
<position>75,-216</position>
<input>
<ID>N_in0</ID>117 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>292</ID>
<type>AA_LABEL</type>
<position>77.5,-211.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>AA_LABEL</type>
<position>77.5,-215.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>294</ID>
<type>AA_LABEL</type>
<position>77.5,-213</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>295</ID>
<type>AA_LABEL</type>
<position>92.5,-199</position>
<gparam>LABEL_TEXT JK TO T</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>297</ID>
<type>BE_JKFF_LOW</type>
<position>108,-213</position>
<input>
<ID>J</ID>119 </input>
<input>
<ID>K</ID>119 </input>
<output>
<ID>Q</ID>121 </output>
<input>
<ID>clock</ID>118 </input>
<output>
<ID>nQ</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>298</ID>
<type>BB_CLOCK</type>
<position>95.5,-213</position>
<output>
<ID>CLK</ID>118 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>299</ID>
<type>AA_TOGGLE</type>
<position>90,-206</position>
<output>
<ID>OUT_0</ID>119 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>301</ID>
<type>GA_LED</type>
<position>115.5,-211</position>
<input>
<ID>N_in0</ID>121 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>302</ID>
<type>GA_LED</type>
<position>116,-215</position>
<input>
<ID>N_in0</ID>122 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>303</ID>
<type>AA_LABEL</type>
<position>118.5,-210.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>304</ID>
<type>AA_LABEL</type>
<position>118.5,-214.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>305</ID>
<type>AA_LABEL</type>
<position>118.5,-212</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>306</ID>
<type>AA_LABEL</type>
<position>49,-204</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>307</ID>
<type>AA_LABEL</type>
<position>90,-203</position>
<gparam>LABEL_TEXT T</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>323</ID>
<type>AA_LABEL</type>
<position>16.5,-227</position>
<gparam>LABEL_TEXT T TO SR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>324</ID>
<type>BE_JKFF_LOW</type>
<position>47.5,-245.5</position>
<input>
<ID>J</ID>138 </input>
<input>
<ID>K</ID>138 </input>
<output>
<ID>Q</ID>132 </output>
<input>
<ID>clock</ID>130 </input>
<output>
<ID>nQ</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>325</ID>
<type>BB_CLOCK</type>
<position>35,-245.5</position>
<output>
<ID>CLK</ID>130 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>327</ID>
<type>GA_LED</type>
<position>55,-243.5</position>
<input>
<ID>N_in0</ID>132 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>328</ID>
<type>GA_LED</type>
<position>55.5,-247.5</position>
<input>
<ID>N_in0</ID>133 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>329</ID>
<type>AA_LABEL</type>
<position>58,-243</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>330</ID>
<type>AA_LABEL</type>
<position>58,-247</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>331</ID>
<type>AA_LABEL</type>
<position>58,-244.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>333</ID>
<type>AA_TOGGLE</type>
<position>15,-240</position>
<output>
<ID>OUT_0</ID>134 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>334</ID>
<type>AA_TOGGLE</type>
<position>15,-248</position>
<output>
<ID>OUT_0</ID>135 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>335</ID>
<type>AA_LABEL</type>
<position>12.5,-239.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>336</ID>
<type>AA_LABEL</type>
<position>12,-247.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>338</ID>
<type>AA_AND2</type>
<position>23,-239</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>134 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>340</ID>
<type>AA_AND2</type>
<position>23.5,-248.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>342</ID>
<type>AE_OR2</type>
<position>33.5,-240</position>
<input>
<ID>IN_0</ID>136 </input>
<input>
<ID>IN_1</ID>137 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>343</ID>
<type>AA_LABEL</type>
<position>78,-227</position>
<gparam>LABEL_TEXT T TO D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>355</ID>
<type>BE_JKFF_LOW</type>
<position>100,-245</position>
<input>
<ID>J</ID>150 </input>
<input>
<ID>K</ID>150 </input>
<output>
<ID>Q</ID>147 </output>
<input>
<ID>clock</ID>145 </input>
<output>
<ID>nQ</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>356</ID>
<type>BB_CLOCK</type>
<position>87.5,-245</position>
<output>
<ID>CLK</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>357</ID>
<type>AA_TOGGLE</type>
<position>73.5,-240</position>
<output>
<ID>OUT_0</ID>149 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>358</ID>
<type>GA_LED</type>
<position>107.5,-243</position>
<input>
<ID>N_in0</ID>147 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>359</ID>
<type>GA_LED</type>
<position>108,-247</position>
<input>
<ID>N_in0</ID>148 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>360</ID>
<type>AA_LABEL</type>
<position>110.5,-242.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>361</ID>
<type>AA_LABEL</type>
<position>110.5,-246.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>362</ID>
<type>AA_LABEL</type>
<position>110.5,-244</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>364</ID>
<type>AI_XOR2</type>
<position>83,-239</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>149 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>365</ID>
<type>AA_LABEL</type>
<position>71.5,-239.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36.5,-25,42,-25</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<intersection>38 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>38,-25,38,-20.5</points>
<intersection>-25 1</intersection>
<intersection>-20.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>30.5,-20.5,38,-20.5</points>
<intersection>30.5 4</intersection>
<intersection>38 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>30.5,-20.5,30.5,-17</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-20.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-15,30.5,-15</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>30.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>30.5,-15,30.5,-15</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-15 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-26,30.5,-26</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<connection>
<GID>6</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-19.5,38,-19.5</points>
<intersection>29.5 3</intersection>
<intersection>38 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>29.5,-24,29.5,-19.5</points>
<intersection>-24 7</intersection>
<intersection>-19.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>38,-19.5,38,-16</points>
<intersection>-19.5 1</intersection>
<intersection>-16 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>36.5,-16,42,-16</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<intersection>38 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>29.5,-24,30.5,-24</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>29.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-14.5,80.5,-14.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-25,92.5,-25</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<intersection>86.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>86.5,-26,86.5,-19</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>-25 1</intersection>
<intersection>-19 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>80.5,-19,86.5,-19</points>
<intersection>80.5 5</intersection>
<intersection>86.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>80.5,-19,80.5,-16.5</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>-19 4</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-16,89.5,-15.5</points>
<intersection>-16 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-16,92.5,-16</points>
<connection>
<GID>23</GID>
<name>N_in0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-15.5,89.5,-15.5</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>88.5 3</intersection>
<intersection>89.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>88.5,-20.5,88.5,-15.5</points>
<intersection>-20.5 4</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>80.5,-20.5,88.5,-20.5</points>
<intersection>80.5 5</intersection>
<intersection>88.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>80.5,-25,80.5,-20.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>-20.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-27,76.5,-26</points>
<intersection>-27 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-26,76.5,-26</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76.5,-27,80.5,-27</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-56.5,43.5,-56.5</points>
<connection>
<GID>54</GID>
<name>N_in0</name></connection>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>39.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>39.5,-56.5,39.5,-52</points>
<intersection>-56.5 1</intersection>
<intersection>-52 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>32,-52,39.5,-52</points>
<intersection>32 4</intersection>
<intersection>39.5 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>32,-52,32,-48.5</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>-52 3</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-51,39.5,-51</points>
<intersection>31 3</intersection>
<intersection>39.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-55.5,31,-51</points>
<intersection>-55.5 7</intersection>
<intersection>-51 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>39.5,-51,39.5,-47.5</points>
<intersection>-51 1</intersection>
<intersection>-47.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>38,-47.5,43.5,-47.5</points>
<connection>
<GID>53</GID>
<name>N_in0</name></connection>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>39.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>31,-55.5,32,-55.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>31 3</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-46.5,32,-46.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<connection>
<GID>63</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-57.5,32,-57.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<connection>
<GID>65</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-56.5,16.5,-47.5</points>
<connection>
<GID>67</GID>
<name>CLK</name></connection>
<intersection>-56.5 2</intersection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-47.5,17,-47.5</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-56.5,18,-56.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-46,14,-45.5</points>
<intersection>-46 2</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14,-45.5,17,-45.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-46,14,-46</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-58.5,14.5,-57</points>
<intersection>-58.5 1</intersection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-58.5,18,-58.5</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10.5,-57,14.5,-57</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>101.5,-56.5,107,-56.5</points>
<connection>
<GID>71</GID>
<name>N_in0</name></connection>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-56.5,103,-52</points>
<intersection>-56.5 1</intersection>
<intersection>-52 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>95.5,-52,103,-52</points>
<intersection>95.5 4</intersection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>95.5,-52,95.5,-48.5</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>-52 3</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94.5,-51,103,-51</points>
<intersection>94.5 3</intersection>
<intersection>103 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>94.5,-55.5,94.5,-51</points>
<intersection>-55.5 7</intersection>
<intersection>-51 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>103,-51,103,-47.5</points>
<intersection>-51 1</intersection>
<intersection>-47.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>101.5,-47.5,107,-47.5</points>
<connection>
<GID>70</GID>
<name>N_in0</name></connection>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>103 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>94.5,-55.5,95.5,-55.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>94.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-46.5,95.5,-46.5</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<connection>
<GID>68</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-57.5,95.5,-57.5</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<connection>
<GID>69</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-56.5,80,-47.5</points>
<connection>
<GID>81</GID>
<name>CLK</name></connection>
<intersection>-56.5 2</intersection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-47.5,80.5,-47.5</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80,-56.5,81.5,-56.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-45.5,80.5,-45.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>70.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>70.5,-48,70.5,-44.5</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>-45.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-58.5,70.5,-52</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70.5,-58.5,81.5,-58.5</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,-71,83,-71</points>
<connection>
<GID>86</GID>
<name>clock</name></connection>
<connection>
<GID>88</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-68,81,-66.5</points>
<intersection>-68 2</intersection>
<intersection>-66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79.5,-66.5,81,-66.5</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81,-68,83,-68</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>89,-68,92,-68</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<connection>
<GID>92</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>89,-71,92.5,-71</points>
<connection>
<GID>86</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>94</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-95,38,-95</points>
<connection>
<GID>111</GID>
<name>clock</name></connection>
<connection>
<GID>113</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-93,35,-90.5</points>
<intersection>-93 1</intersection>
<intersection>-90.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-93,38,-93</points>
<connection>
<GID>111</GID>
<name>J</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-90.5,35,-90.5</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-99,35.5,-97</points>
<intersection>-99 2</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-97,38,-97</points>
<connection>
<GID>111</GID>
<name>K</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-99,35.5,-99</points>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-93,47.5,-93</points>
<connection>
<GID>119</GID>
<name>N_in0</name></connection>
<connection>
<GID>111</GID>
<name>Q</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-97,47.5,-97</points>
<connection>
<GID>121</GID>
<name>N_in0</name></connection>
<connection>
<GID>111</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-96,88.5,-96</points>
<connection>
<GID>153</GID>
<name>CLK</name></connection>
<connection>
<GID>152</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94.5,-94,98,-94</points>
<connection>
<GID>156</GID>
<name>N_in0</name></connection>
<connection>
<GID>152</GID>
<name>Q</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94.5,-98,98,-98</points>
<connection>
<GID>157</GID>
<name>N_in0</name></connection>
<connection>
<GID>152</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-98.5,76,-90</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<intersection>-98.5 3</intersection>
<intersection>-93.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-93.5,88.5,-93.5</points>
<intersection>76 0</intersection>
<intersection>88.5 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>76,-98.5,88.5,-98.5</points>
<intersection>76 0</intersection>
<intersection>88.5 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>88.5,-94,88.5,-93.5</points>
<connection>
<GID>152</GID>
<name>J</name></connection>
<intersection>-93.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>88.5,-98.5,88.5,-98</points>
<connection>
<GID>152</GID>
<name>K</name></connection>
<intersection>-98.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-125.5,40.5,-123.5</points>
<intersection>-125.5 2</intersection>
<intersection>-123.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-123.5,40.5,-123.5</points>
<connection>
<GID>165</GID>
<name>OUTINV_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-125.5,50,-125.5</points>
<connection>
<GID>169</GID>
<name>N_in0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-136.5,32.5,-136.5</points>
<connection>
<GID>173</GID>
<name>CLK</name></connection>
<intersection>32.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>32.5,-136.5,32.5,-123.5</points>
<connection>
<GID>165</GID>
<name>clock</name></connection>
<intersection>-136.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-116,18.5,-115</points>
<connection>
<GID>171</GID>
<name>OUT_0</name></connection>
<connection>
<GID>177</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-121,18.5,-120</points>
<connection>
<GID>177</GID>
<name>OUT_0</name></connection>
<connection>
<GID>179</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-121,20.5,-116.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-116.5,47,-116.5</points>
<intersection>20.5 0</intersection>
<intersection>47 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>47,-121,47,-116.5</points>
<intersection>-121 4</intersection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>38.5,-121,51,-121</points>
<connection>
<GID>167</GID>
<name>N_in0</name></connection>
<intersection>38.5 5</intersection>
<intersection>47 2</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>38.5,-121,38.5,-120.5</points>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<intersection>-121 4</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-127.5,14.5,-115</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<connection>
<GID>175</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-127.5,16.5,-127</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>-127 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-127,19.5,-127</points>
<connection>
<GID>179</GID>
<name>OUT</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-133.5,24,-120.5</points>
<intersection>-133.5 2</intersection>
<intersection>-120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-120.5,32.5,-120.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-133.5,24,-133.5</points>
<connection>
<GID>181</GID>
<name>OUT</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99.5,-151,105,-151</points>
<connection>
<GID>190</GID>
<name>N_in0</name></connection>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-151,101,-146.5</points>
<intersection>-151 1</intersection>
<intersection>-146.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>93.5,-146.5,101,-146.5</points>
<intersection>93.5 4</intersection>
<intersection>101 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93.5,-146.5,93.5,-143</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<intersection>-146.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-137.5,100.5,-137.5</points>
<intersection>59 8</intersection>
<intersection>100.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>100.5,-147,100.5,-137.5</points>
<intersection>-147 7</intersection>
<intersection>-142 6</intersection>
<intersection>-137.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>99.5,-142,105,-142</points>
<connection>
<GID>189</GID>
<name>N_in0</name></connection>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<intersection>100.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>93.5,-147,100.5,-147</points>
<intersection>93.5 9</intersection>
<intersection>100.5 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>59,-142,59,-137.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>-137.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>93.5,-150,93.5,-147</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>-147 7</intersection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-141,93.5,-141</points>
<connection>
<GID>196</GID>
<name>OUT</name></connection>
<connection>
<GID>187</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-152,93.5,-152</points>
<connection>
<GID>197</GID>
<name>OUT</name></connection>
<connection>
<GID>188</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-151,78,-142</points>
<connection>
<GID>198</GID>
<name>CLK</name></connection>
<intersection>-151 2</intersection>
<intersection>-142 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-142,78.5,-142</points>
<connection>
<GID>196</GID>
<name>IN_1</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-151,79.5,-151</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65.5,-140,78.5,-140</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>65.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>65.5,-154.5,65.5,-140</points>
<intersection>-154.5 5</intersection>
<intersection>-142.5 6</intersection>
<intersection>-140 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>54,-154.5,65.5,-154.5</points>
<connection>
<GID>204</GID>
<name>OUT</name></connection>
<intersection>65.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>65.5,-142.5,68.5,-142.5</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>65.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-153,68.5,-146.5</points>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection>
<intersection>-153 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-153,79.5,-153</points>
<connection>
<GID>197</GID>
<name>IN_1</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-142,57,-141</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-148.5,55,-148</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>-148 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>55,-148,58,-148</points>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-142,52.5,-136</points>
<connection>
<GID>200</GID>
<name>OUT_0</name></connection>
<intersection>-142 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>53,-148.5,53,-142</points>
<connection>
<GID>204</GID>
<name>IN_1</name></connection>
<intersection>-142 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>52.5,-142,53,-142</points>
<intersection>52.5 0</intersection>
<intersection>53 1</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>56.5,-137,56.5,-136</points>
<connection>
<GID>201</GID>
<name>OUT_0</name></connection>
<intersection>-137 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>56.5,-137,57,-137</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>56.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,-185,42,-185</points>
<intersection>18.5 3</intersection>
<intersection>42 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18.5,-185,18.5,-181.5</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<intersection>-185 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>42,-185,42,-174</points>
<intersection>-185 1</intersection>
<intersection>-174 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>39,-174,46,-174</points>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection>
<connection>
<GID>217</GID>
<name>N_in0</name></connection>
<intersection>42 4</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15.5,-167,43.5,-167</points>
<intersection>15.5 4</intersection>
<intersection>43.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43.5,-177,43.5,-167</points>
<intersection>-177 6</intersection>
<intersection>-167 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>15.5,-170.5,15.5,-167</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>-167 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>39,-177,46,-177</points>
<connection>
<GID>209</GID>
<name>OUTINV_0</name></connection>
<intersection>43.5 3</intersection>
<intersection>46 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>46,-177.5,46,-177</points>
<connection>
<GID>219</GID>
<name>N_in0</name></connection>
<intersection>-177 6</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-190,31,-177</points>
<intersection>-190 1</intersection>
<intersection>-177 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-190,31,-190</points>
<connection>
<GID>215</GID>
<name>CLK</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-177,33,-177</points>
<connection>
<GID>209</GID>
<name>clock</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-172.5,15.5,-172.5</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<connection>
<GID>211</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-179.5,14,-179.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<connection>
<GID>213</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-179.5,18.5,-179.5</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<connection>
<GID>225</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-173.5,22.5,-171.5</points>
<intersection>-173.5 2</intersection>
<intersection>-171.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-171.5,22.5,-171.5</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-173.5,24.5,-173.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-180.5,24.5,-175.5</points>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<connection>
<GID>225</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-174.5,31,-174</points>
<intersection>-174.5 2</intersection>
<intersection>-174 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-174,33,-174</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-174.5,31,-174.5</points>
<connection>
<GID>227</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-168.5,91,-168.5</points>
<intersection>72 3</intersection>
<intersection>91 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>72,-171.5,72,-168.5</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>-168.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>91,-174.5,91,-168.5</points>
<intersection>-174.5 6</intersection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>89,-174.5,92.5,-174.5</points>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection>
<connection>
<GID>241</GID>
<name>N_in0</name></connection>
<intersection>91 4</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-178,90.5,-177.5</points>
<intersection>-178 1</intersection>
<intersection>-177.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90.5,-178,92.5,-178</points>
<connection>
<GID>242</GID>
<name>N_in0</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89,-177.5,90.5,-177.5</points>
<connection>
<GID>240</GID>
<name>OUTINV_0</name></connection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-183,82,-177.5</points>
<intersection>-183 1</intersection>
<intersection>-177.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,-183,82,-183</points>
<connection>
<GID>246</GID>
<name>CLK</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-177.5,83,-177.5</points>
<connection>
<GID>240</GID>
<name>clock</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-173.5,70,-173</points>
<intersection>-173.5 1</intersection>
<intersection>-173 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-173.5,72,-173.5</points>
<connection>
<GID>249</GID>
<name>IN_1</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68.5,-173,70,-173</points>
<connection>
<GID>247</GID>
<name>OUT_0</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-174.5,80.5,-172.5</points>
<intersection>-174.5 1</intersection>
<intersection>-172.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-174.5,83,-174.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-172.5,80.5,-172.5</points>
<connection>
<GID>249</GID>
<name>OUT</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-213.5,22,-212</points>
<intersection>-213.5 1</intersection>
<intersection>-212 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-213.5,26.5,-213.5</points>
<connection>
<GID>253</GID>
<name>J</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-212,22,-212</points>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-220,22.5,-217.5</points>
<intersection>-220 2</intersection>
<intersection>-217.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-217.5,26.5,-217.5</points>
<connection>
<GID>253</GID>
<name>K</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-220,22.5,-220</points>
<connection>
<GID>257</GID>
<name>OUT_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-215.5,26.5,-215.5</points>
<connection>
<GID>253</GID>
<name>clock</name></connection>
<connection>
<GID>259</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-213.5,34,-213</points>
<intersection>-213.5 2</intersection>
<intersection>-213 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-213,35.5,-213</points>
<connection>
<GID>261</GID>
<name>N_in0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-213.5,34,-213.5</points>
<connection>
<GID>253</GID>
<name>Q</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32.5,-217.5,35.5,-217.5</points>
<connection>
<GID>263</GID>
<name>N_in0</name></connection>
<connection>
<GID>253</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-214,64,-214</points>
<connection>
<GID>287</GID>
<name>CLK</name></connection>
<connection>
<GID>286</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-212.5,49,-209</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<connection>
<GID>288</GID>
<name>OUT_0</name></connection>
<intersection>-211 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-211,64,-211</points>
<intersection>49 0</intersection>
<intersection>64 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>64,-212,64,-211</points>
<connection>
<GID>286</GID>
<name>J</name></connection>
<intersection>-211 1</intersection></vsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-217,49,-216.5</points>
<connection>
<GID>289</GID>
<name>OUT_0</name></connection>
<intersection>-217 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-217,64,-217</points>
<intersection>49 0</intersection>
<intersection>64 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>64,-217,64,-216</points>
<connection>
<GID>286</GID>
<name>K</name></connection>
<intersection>-217 1</intersection></vsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-212,73.5,-212</points>
<connection>
<GID>286</GID>
<name>Q</name></connection>
<connection>
<GID>290</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-216,74,-216</points>
<connection>
<GID>286</GID>
<name>nQ</name></connection>
<connection>
<GID>291</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99.5,-213,105,-213</points>
<connection>
<GID>298</GID>
<name>CLK</name></connection>
<connection>
<GID>297</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-215,90,-208</points>
<connection>
<GID>299</GID>
<name>OUT_0</name></connection>
<intersection>-215 7</intersection>
<intersection>-210 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>90,-215,105,-215</points>
<connection>
<GID>297</GID>
<name>K</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>90,-210,105,-210</points>
<intersection>90 0</intersection>
<intersection>105 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>105,-211,105,-210</points>
<connection>
<GID>297</GID>
<name>J</name></connection>
<intersection>-210 8</intersection></vsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,-211,114.5,-211</points>
<connection>
<GID>301</GID>
<name>N_in0</name></connection>
<connection>
<GID>297</GID>
<name>Q</name></connection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,-215,115,-215</points>
<connection>
<GID>302</GID>
<name>N_in0</name></connection>
<connection>
<GID>297</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-245.5,44.5,-245.5</points>
<connection>
<GID>325</GID>
<name>CLK</name></connection>
<connection>
<GID>324</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-252.5,53,-252.5</points>
<intersection>20.5 4</intersection>
<intersection>53 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20.5,-252.5,20.5,-249.5</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<intersection>-252.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>53,-252.5,53,-243.5</points>
<intersection>-252.5 1</intersection>
<intersection>-243.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>50.5,-243.5,54,-243.5</points>
<connection>
<GID>324</GID>
<name>Q</name></connection>
<connection>
<GID>327</GID>
<name>N_in0</name></connection>
<intersection>53 5</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,-236,52,-236</points>
<intersection>20 4</intersection>
<intersection>52 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,-238,20,-236</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>-236 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>52,-247.5,52,-236</points>
<intersection>-247.5 7</intersection>
<intersection>-236 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>50.5,-247.5,54.5,-247.5</points>
<connection>
<GID>324</GID>
<name>nQ</name></connection>
<connection>
<GID>328</GID>
<name>N_in0</name></connection>
<intersection>52 5</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-240,20,-240</points>
<connection>
<GID>333</GID>
<name>OUT_0</name></connection>
<connection>
<GID>338</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-248,18.5,-247.5</points>
<intersection>-248 1</intersection>
<intersection>-247.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-248,18.5,-248</points>
<connection>
<GID>334</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-247.5,20.5,-247.5</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-239,30.5,-239</points>
<connection>
<GID>338</GID>
<name>OUT</name></connection>
<connection>
<GID>342</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-248.5,28.5,-241</points>
<intersection>-248.5 1</intersection>
<intersection>-241 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-248.5,28.5,-248.5</points>
<connection>
<GID>340</GID>
<name>OUT</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-241,30.5,-241</points>
<connection>
<GID>342</GID>
<name>IN_1</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-242.5,40.5,-240</points>
<intersection>-242.5 1</intersection>
<intersection>-240 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-242.5,44.5,-242.5</points>
<intersection>31 3</intersection>
<intersection>40.5 0</intersection>
<intersection>44.5 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-240,40.5,-240</points>
<connection>
<GID>342</GID>
<name>OUT</name></connection>
<intersection>40.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-248,31,-242.5</points>
<intersection>-248 4</intersection>
<intersection>-242.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>31,-248,44.5,-248</points>
<intersection>31 3</intersection>
<intersection>44.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>44.5,-248,44.5,-247.5</points>
<connection>
<GID>324</GID>
<name>K</name></connection>
<intersection>-248 4</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>44.5,-243.5,44.5,-242.5</points>
<connection>
<GID>324</GID>
<name>J</name></connection>
<intersection>-242.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91.5,-245,97,-245</points>
<connection>
<GID>356</GID>
<name>CLK</name></connection>
<connection>
<GID>355</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>77.5,-235.5,104,-235.5</points>
<intersection>77.5 4</intersection>
<intersection>104 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>77.5,-238,77.5,-235.5</points>
<intersection>-238 7</intersection>
<intersection>-235.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>104,-243,104,-235.5</points>
<intersection>-243 8</intersection>
<intersection>-235.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>77.5,-238,80,-238</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>77.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>103,-243,106.5,-243</points>
<connection>
<GID>355</GID>
<name>Q</name></connection>
<connection>
<GID>358</GID>
<name>N_in0</name></connection>
<intersection>104 5</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-247,107,-247</points>
<connection>
<GID>359</GID>
<name>N_in0</name></connection>
<connection>
<GID>355</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75.5,-240,80,-240</points>
<connection>
<GID>364</GID>
<name>IN_1</name></connection>
<connection>
<GID>357</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-242,91.5,-239</points>
<intersection>-242 1</intersection>
<intersection>-239 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-242,97,-242</points>
<intersection>82.5 3</intersection>
<intersection>91.5 0</intersection>
<intersection>97 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86,-239,91.5,-239</points>
<connection>
<GID>364</GID>
<name>OUT</name></connection>
<intersection>91.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>82.5,-249,82.5,-242</points>
<intersection>-249 4</intersection>
<intersection>-242 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>82.5,-249,97,-249</points>
<intersection>82.5 3</intersection>
<intersection>97 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>97,-243,97,-242</points>
<connection>
<GID>355</GID>
<name>J</name></connection>
<intersection>-242 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>97,-249,97,-247</points>
<connection>
<GID>355</GID>
<name>K</name></connection>
<intersection>-249 4</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>